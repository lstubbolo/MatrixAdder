library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.std_logic_textio.all;
use IEEE.std_logic_arith.all;
use IEEE.numeric_bit.all;
use IEEE.numeric_std.all;
use IEEE.std_logic_signed.all;
--use IEEE.std_logic_unsigned.all;

entity matrix_0_v1_0_S00_AXI is
	generic (
		C_S_AXI_DATA_WIDTH	: integer	:= 32;
		C_S_AXI_ADDR_WIDTH	: integer	:= 11
	);
	port (
		-- Global Clock Signal
		S_AXI_ACLK    : in std_logic;
		S_AXI_ARESETN : in std_logic;
		
		-- Write address (issued by master, acceped by Slave)
		S_AXI_AWADDR	: in std_logic_vector(C_S_AXI_ADDR_WIDTH-1 downto 0);
		
		S_AXI_AWPROT  : in std_logic_vector(2 downto 0);
		S_AXI_AWVALID : in std_logic;
		S_AXI_AWREADY : out std_logic;
		S_AXI_WDATA	  : in std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
		S_AXI_WSTRB	  : in std_logic_vector((C_S_AXI_DATA_WIDTH/8)-1 downto 0);
		S_AXI_WVALID  : in std_logic;
		S_AXI_WREADY  : out std_logic;
		S_AXI_BRESP   : out std_logic_vector(1 downto 0);
		S_AXI_BVALID  : out std_logic;
		S_AXI_BREADY  : in std_logic;
		S_AXI_ARADDR  : in std_logic_vector(C_S_AXI_ADDR_WIDTH-1 downto 0);
		S_AXI_ARPROT  : in std_logic_vector(2 downto 0);
		S_AXI_ARVALID : in std_logic;
		S_AXI_ARREADY : out std_logic;
		S_AXI_RDATA	  : out std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
		S_AXI_RRESP	  : out std_logic_vector(1 downto 0);
		S_AXI_RVALID  : out std_logic;
		S_AXI_RREADY  : in std_logic
	);
end matrix_0_v1_0_S00_AXI;

--  = # = # = # = # = # = # = # = # = # = # = # = # = # = # = # = # = # = # = # = # = # = # = # = # = # = # = # = #

--                        A R C H I T E C T U R E    S T A T E M E N T    

architecture arch_imp of matrix_0_v1_0_S00_AXI is

	-- AXI4LITE signals
	signal axi_awaddr	: std_logic_vector(C_S_AXI_ADDR_WIDTH-1 downto 0);
	signal axi_awready	: std_logic;
	signal axi_wready	: std_logic;
	signal axi_bresp	: std_logic_vector(1 downto 0);
	signal axi_bvalid	: std_logic;
	signal axi_araddr	: std_logic_vector(C_S_AXI_ADDR_WIDTH-1 downto 0);
	signal axi_arready	: std_logic;
	signal axi_rdata	: std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
	signal axi_rresp	: std_logic_vector(1 downto 0);
	signal axi_rvalid	: std_logic;

	constant ADDR_LSB  : integer := (C_S_AXI_DATA_WIDTH/32)+ 1;
	constant OPT_MEM_ADDR_BITS : integer := 8;

    constant N          : integer := 16;





--  = # = # = # = # = # = # = # = # = # = # = # = # = # = # = # = # = # = # = # = # = # = # = # = # = # = # = # = #

            --  S L A V E    R E G I S T E R    S I G N A L    D E C L A R A T I O N	
	
	-- 
	signal slv_reg0    :std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0) := (others => '1');
    signal slv_reg256  :std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0) := (others => '1');
	
    signal 

            --  Registers used for A input: 0 - 127

--  0              1              2              3              4              5              6              7
	         	   slv_reg1,	  slv_reg2,	     slv_reg3,	    slv_reg4,	   slv_reg5,	  slv_reg6,	     slv_reg7,	
	slv_reg8,	   slv_reg9,	  slv_reg10,	 slv_reg11,	    slv_reg12,	   slv_reg13,	  slv_reg14,	 slv_reg15,	
	slv_reg16,	   slv_reg17,	  slv_reg18,	 slv_reg19,	    slv_reg20,	   slv_reg21,	  slv_reg22,	 slv_reg23,	
	slv_reg24,	   slv_reg25,	  slv_reg26,	 slv_reg27,	    slv_reg28,	   slv_reg29,	  slv_reg30,	 slv_reg31,	
	slv_reg32,	   slv_reg33,	  slv_reg34,	 slv_reg35,	    slv_reg36,	   slv_reg37,	  slv_reg38,	 slv_reg39,	
	slv_reg40,	   slv_reg41,	  slv_reg42,	 slv_reg43,	    slv_reg44,	   slv_reg45,	  slv_reg46,	 slv_reg47,	
	slv_reg48,	   slv_reg49,	  slv_reg50,	 slv_reg51,	    slv_reg52,	   slv_reg53,	  slv_reg54,	 slv_reg55,	
	slv_reg56,	   slv_reg57,	  slv_reg58,	 slv_reg59,	    slv_reg60,	   slv_reg61,	  slv_reg62,	 slv_reg63,	
	slv_reg64,	   slv_reg65,	  slv_reg66,	 slv_reg67,	    slv_reg68,	   slv_reg69,	  slv_reg70,	 slv_reg71,	
	slv_reg72,	   slv_reg73,	  slv_reg74,	 slv_reg75,	    slv_reg76,	   slv_reg77,	  slv_reg78,	 slv_reg79,	
	slv_reg80,	   slv_reg81,	  slv_reg82,	 slv_reg83,	    slv_reg84,	   slv_reg85,	  slv_reg86,	 slv_reg87,	
	slv_reg88,	   slv_reg89,	  slv_reg90,	 slv_reg91,	    slv_reg92,	   slv_reg93,	  slv_reg94,	 slv_reg95,	
	slv_reg96,	   slv_reg97,	  slv_reg98,	 slv_reg99,	    slv_reg100,	   slv_reg101,	  slv_reg102,	 slv_reg103,	
	slv_reg104,	   slv_reg105,	  slv_reg106,	 slv_reg107,	slv_reg108,	   slv_reg109,	  slv_reg110,	 slv_reg111,	
	slv_reg112,	   slv_reg113,	  slv_reg114,	 slv_reg115,	slv_reg116,	   slv_reg117,	  slv_reg118,	 slv_reg119,	
	slv_reg120,	   slv_reg121,	  slv_reg122,	 slv_reg123,	slv_reg124,	   slv_reg125,	  slv_reg126,	 slv_reg127,

--  = # = # = # = # = # = # = # = # = # = # = # = # = # = # = # = # = # = # = # = # = # = # = # = # = # = # = # = #
            
            --  Registers used for B input: 128 - 255
            
--  0              1              2              3              4              5              6              7
    slv_reg128,	   slv_reg129,    slv_reg130,	 slv_reg131,	slv_reg132,    slv_reg133,	  slv_reg134,	 slv_reg135,	
    slv_reg136,    slv_reg137,    slv_reg138,    slv_reg139,    slv_reg140,    slv_reg141,    slv_reg142,    slv_reg143,    
    slv_reg144,    slv_reg145,    slv_reg146,    slv_reg147,    slv_reg148,    slv_reg149,    slv_reg150,    slv_reg151,    
    slv_reg152,    slv_reg153,    slv_reg154,    slv_reg155,    slv_reg156,    slv_reg157,    slv_reg158,    slv_reg159,    
    slv_reg160,    slv_reg161,    slv_reg162,    slv_reg163,    slv_reg164,    slv_reg165,    slv_reg166,    slv_reg167,    
    slv_reg168,    slv_reg169,    slv_reg170,    slv_reg171,    slv_reg172,    slv_reg173,    slv_reg174,    slv_reg175,    
    slv_reg176,    slv_reg177,    slv_reg178,    slv_reg179,    slv_reg180,    slv_reg181,    slv_reg182,    slv_reg183,    
    slv_reg184,    slv_reg185,    slv_reg186,    slv_reg187,    slv_reg188,    slv_reg189,    slv_reg190,    slv_reg191,    
    slv_reg192,    slv_reg193,    slv_reg194,    slv_reg195,    slv_reg196,    slv_reg197,    slv_reg198,    slv_reg199,    
    slv_reg200,    slv_reg201,    slv_reg202,    slv_reg203,    slv_reg204,    slv_reg205,    slv_reg206,    slv_reg207,    
    slv_reg208,    slv_reg209,    slv_reg210,    slv_reg211,    slv_reg212,    slv_reg213,    slv_reg214,    slv_reg215,    
    slv_reg216,    slv_reg217,    slv_reg218,    slv_reg219,    slv_reg220,    slv_reg221,    slv_reg222,    slv_reg223,    
    slv_reg224,    slv_reg225,    slv_reg226,    slv_reg227,    slv_reg228,    slv_reg229,    slv_reg230,    slv_reg231,    
    slv_reg232,    slv_reg233,    slv_reg234,    slv_reg235,    slv_reg236,    slv_reg237,    slv_reg238,    slv_reg239,    
    slv_reg240,    slv_reg241,    slv_reg242,    slv_reg243,    slv_reg244,    slv_reg245,    slv_reg246,    slv_reg247,    
    slv_reg248,    slv_reg249,    slv_reg250,    slv_reg251,    slv_reg252,    slv_reg253,    slv_reg254,    slv_reg255,	

--  = # = # = # = # = # = # = # = # = # = # = # = # = # = # = # = # = # = # = # = # = # = # = # = # = # = # = # = #
            
            --  Registers used for C Output (256 - 511)
            
--  0              1              2              3              4              5              6              7
	               slv_reg257,     slv_reg258,   slv_reg259,    slv_reg260,    slv_reg261,    slv_reg262,    slv_reg263, 
    slv_reg264,    slv_reg265,     slv_reg266,   slv_reg267,    slv_reg268,    slv_reg269,    slv_reg270,    slv_reg271, 
    slv_reg272,    slv_reg273,     slv_reg274,   slv_reg275,    slv_reg276,    slv_reg277,    slv_reg278,    slv_reg279, 
    slv_reg280,    slv_reg281,     slv_reg282,   slv_reg283,    slv_reg284,    slv_reg285,    slv_reg286,    slv_reg287, 
    slv_reg288,    slv_reg289,     slv_reg290,   slv_reg291,    slv_reg292,    slv_reg293,    slv_reg294,    slv_reg295, 
    slv_reg296,    slv_reg297,     slv_reg298,   slv_reg299,    slv_reg300,    slv_reg301,    slv_reg302,    slv_reg303, 
    slv_reg304,    slv_reg305,     slv_reg306,   slv_reg307,    slv_reg308,    slv_reg309,    slv_reg310,    slv_reg311, 
    slv_reg312,    slv_reg313,     slv_reg314,   slv_reg315,    slv_reg316,    slv_reg317,    slv_reg318,    slv_reg319, 
    slv_reg320,    slv_reg321,     slv_reg322,   slv_reg323,    slv_reg324,    slv_reg325,    slv_reg326,    slv_reg327, 
    slv_reg328,    slv_reg329,     slv_reg330,   slv_reg331,    slv_reg332,    slv_reg333,    slv_reg334,    slv_reg335, 
    slv_reg336,    slv_reg337,     slv_reg338,   slv_reg339,    slv_reg340,    slv_reg341,    slv_reg342,    slv_reg343, 
    slv_reg344,    slv_reg345,     slv_reg346,   slv_reg347,    slv_reg348,    slv_reg349,    slv_reg350,    slv_reg351, 
    slv_reg352,    slv_reg353,     slv_reg354,   slv_reg355,    slv_reg356,    slv_reg357,    slv_reg358,    slv_reg359, 
    slv_reg360,    slv_reg361,     slv_reg362,   slv_reg363,    slv_reg364,    slv_reg365,    slv_reg366,    slv_reg367, 
    slv_reg368,    slv_reg369,     slv_reg370,   slv_reg371,    slv_reg372,    slv_reg373,    slv_reg374,    slv_reg375, 
    slv_reg376,    slv_reg377,     slv_reg378,   slv_reg379,    slv_reg380,    slv_reg381,    slv_reg382,    slv_reg383, 
    slv_reg384,    slv_reg385,     slv_reg386,   slv_reg387,    slv_reg388,    slv_reg389,    slv_reg390,    slv_reg391, 
    slv_reg392,    slv_reg393,     slv_reg394,   slv_reg395,    slv_reg396,    slv_reg397,    slv_reg398,    slv_reg399, 
    slv_reg400,    slv_reg401,     slv_reg402,   slv_reg403,    slv_reg404,    slv_reg405,    slv_reg406,    slv_reg407, 
    slv_reg408,    slv_reg409,     slv_reg410,   slv_reg411,    slv_reg412,    slv_reg413,    slv_reg414,    slv_reg415, 
    slv_reg416,    slv_reg417,     slv_reg418,   slv_reg419,    slv_reg420,    slv_reg421,    slv_reg422,    slv_reg423, 
    slv_reg424,    slv_reg425,     slv_reg426,   slv_reg427,    slv_reg428,    slv_reg429,    slv_reg430,    slv_reg431, 
    slv_reg432,    slv_reg433,     slv_reg434,   slv_reg435,    slv_reg436,    slv_reg437,    slv_reg438,    slv_reg439, 
    slv_reg440,    slv_reg441,     slv_reg442,   slv_reg443,    slv_reg444,    slv_reg445,    slv_reg446,    slv_reg447, 
    slv_reg448,    slv_reg449,     slv_reg450,   slv_reg451,    slv_reg452,    slv_reg453,    slv_reg454,    slv_reg455, 
    slv_reg456,    slv_reg457,     slv_reg458,   slv_reg459,    slv_reg460,    slv_reg461,    slv_reg462,    slv_reg463, 
    slv_reg464,    slv_reg465,     slv_reg466,   slv_reg467,    slv_reg468,    slv_reg469,    slv_reg470,    slv_reg471, 
    slv_reg472,    slv_reg473,     slv_reg474,   slv_reg475,    slv_reg476,    slv_reg477,    slv_reg478,    slv_reg479, 
    slv_reg480,    slv_reg481,     slv_reg482,   slv_reg483,    slv_reg484,    slv_reg485,    slv_reg486,    slv_reg487, 
    slv_reg488,    slv_reg489,     slv_reg490,   slv_reg491,    slv_reg492,    slv_reg493,    slv_reg494,    slv_reg495, 
    slv_reg496,    slv_reg497,     slv_reg498,   slv_reg499,    slv_reg500,    slv_reg501,    slv_reg502,    slv_reg503, 
    slv_reg504,    slv_reg505,     slv_reg506,   slv_reg507,    slv_reg508,    slv_reg509,    slv_reg510,    slv_reg511
    	
:std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);


	signal slv_reg_rden    : std_logic;
	signal slv_reg_wren    : std_logic;
	signal reg_data_out    : std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
	signal byte_index      : integer;
	signal aw_en           : std_logic;


--  = # = # = # = # = # = # = # = # = # = # = # = # = # = # = # = # = # = # = # = # = # = # = # = # = # = # = # = #

--                        U S E R    S I G N A L S  /  C O M P O N E N T S


--  Start massive copy / paste here -> Ends at ctrl + F (***NOTE)

--  output signals

signal	out_0_0,	out_0_1,	out_0_2,	out_0_3,	out_0_4,	out_0_5,	out_0_6,	out_0_7,	

        out_1_0,    out_1_1,    out_1_2,    out_1_3,    out_1_4,    out_1_5,    out_1_6,    out_1_7,    

        out_2_0,    out_2_1,    out_2_2,    out_2_3,    out_2_4,    out_2_5,    out_2_6,    out_2_7,    

        out_3_0,    out_3_1,    out_3_2,    out_3_3,    out_3_4,    out_3_5,    out_3_6,    out_3_7,    

        out_4_0,    out_4_1,    out_4_2,    out_4_3,    out_4_4,    out_4_5,    out_4_6,    out_4_7,    

        out_5_0,    out_5_1,    out_5_2,    out_5_3,    out_5_4,    out_5_5,    out_5_6,    out_5_7,    

        out_6_0,    out_6_1,    out_6_2,    out_6_3,    out_6_4,    out_6_5,    out_6_6,    out_6_7,    

        out_7_0,    out_7_1,    out_7_2,    out_7_3,    out_7_4,    out_7_5,    out_7_6,    out_7_7    

: STD_LOGIC_VECTOR(31 downto 0);  



    
    
    
--  = # = # = # = # = # = # = # = # = # = # = # = # = # = # = # = # = # = # = # = # = # = # = # = # = # = # = # = #

--                                B E G I N    S T A T E M E N T


begin



--  = # = # = # = # = # = # = # = # = # = # = # = # = # = # = # = # = # = # = # = # = # = # = # = # = # = # = # = # 
--  = # = # = # = # = # = # = # = # = # = # = # = # = # = # = # = # = # = # = # = # = # = # = # = # = # = # = # = #


       --                                          U S E R    L O G I C   

    
--  = # = # = # = # = # = # = # = # = # = # = # = # = # = # = # = # = # = # = # = # = # = # = # = # = # = # = # = # 
--  = # = # = # = # = # = # = # = # = # = # = # = # = # = # = # = # = # = # = # = # = # = # = # = # = # = # = # = #








--  = # = # = # = # = # = # = # = # = # = # = # = # = # = # = # = # = # = # = # = # = # = # = # = # = # = # = # = # 
--  = # = # = # = # = # = # = # = # = # = # = # = # = # = # = # = # = # = # = # = # = # = # = # = # = # = # = # = #


       --                                   O U T P U T   C A L C U L A T I O N S


--  = # = # = # = # = # = # = # = # = # = # = # = # = # = # = # = # = # = # = # = # = # = # = # = # = # = # = # = # 
--  = # = # = # = # = # = # = # = # = # = # = # = # = # = # = # = # = # = # = # = # = # = # = # = # = # = # = # = #



out_0_0 <= 		   slv_reg0(15 downto 0) * slv_reg128(15 downto 0)	 + slv_reg1(15 downto 0) * slv_reg136(15 downto 0)
				 + slv_reg2(15 downto 0) * slv_reg144(15 downto 0)	 + slv_reg3(15 downto 0) * slv_reg152(15 downto 0)
				 + slv_reg4(15 downto 0) * slv_reg160(15 downto 0)	 + slv_reg5(15 downto 0) * slv_reg168(15 downto 0)
				 + slv_reg6(15 downto 0) * slv_reg176(15 downto 0)	 + slv_reg7(15 downto 0) * slv_reg184(15 downto 0);
out_0_1 <= 		   slv_reg0(15 downto 0) * slv_reg129(15 downto 0)	 + slv_reg1(15 downto 0) * slv_reg137(15 downto 0)
				 + slv_reg2(15 downto 0) * slv_reg145(15 downto 0)	 + slv_reg3(15 downto 0) * slv_reg153(15 downto 0)
				 + slv_reg4(15 downto 0) * slv_reg161(15 downto 0)	 + slv_reg5(15 downto 0) * slv_reg169(15 downto 0)
				 + slv_reg6(15 downto 0) * slv_reg177(15 downto 0)	 + slv_reg7(15 downto 0) * slv_reg185(15 downto 0);
out_0_2 <= 		   slv_reg0(15 downto 0) * slv_reg130(15 downto 0)	 + slv_reg1(15 downto 0) * slv_reg138(15 downto 0)
				 + slv_reg2(15 downto 0) * slv_reg146(15 downto 0)	 + slv_reg3(15 downto 0) * slv_reg154(15 downto 0)
				 + slv_reg4(15 downto 0) * slv_reg162(15 downto 0)	 + slv_reg5(15 downto 0) * slv_reg170(15 downto 0)
				 + slv_reg6(15 downto 0) * slv_reg178(15 downto 0)	 + slv_reg7(15 downto 0) * slv_reg186(15 downto 0);
out_0_3 <= 		   slv_reg0(15 downto 0) * slv_reg131(15 downto 0)	 + slv_reg1(15 downto 0) * slv_reg139(15 downto 0)
				 + slv_reg2(15 downto 0) * slv_reg147(15 downto 0)	 + slv_reg3(15 downto 0) * slv_reg155(15 downto 0)
				 + slv_reg4(15 downto 0) * slv_reg163(15 downto 0)	 + slv_reg5(15 downto 0) * slv_reg171(15 downto 0)
				 + slv_reg6(15 downto 0) * slv_reg179(15 downto 0)	 + slv_reg7(15 downto 0) * slv_reg187(15 downto 0);
out_0_4 <= 		   slv_reg0(15 downto 0) * slv_reg132(15 downto 0)	 + slv_reg1(15 downto 0) * slv_reg140(15 downto 0)
				 + slv_reg2(15 downto 0) * slv_reg148(15 downto 0)	 + slv_reg3(15 downto 0) * slv_reg156(15 downto 0)
				 + slv_reg4(15 downto 0) * slv_reg164(15 downto 0)	 + slv_reg5(15 downto 0) * slv_reg172(15 downto 0)
				 + slv_reg6(15 downto 0) * slv_reg180(15 downto 0)	 + slv_reg7(15 downto 0) * slv_reg188(15 downto 0);
out_0_5 <= 		   slv_reg0(15 downto 0) * slv_reg133(15 downto 0)	 + slv_reg1(15 downto 0) * slv_reg141(15 downto 0)
				 + slv_reg2(15 downto 0) * slv_reg149(15 downto 0)	 + slv_reg3(15 downto 0) * slv_reg157(15 downto 0)
				 + slv_reg4(15 downto 0) * slv_reg165(15 downto 0)	 + slv_reg5(15 downto 0) * slv_reg173(15 downto 0)
				 + slv_reg6(15 downto 0) * slv_reg181(15 downto 0)	 + slv_reg7(15 downto 0) * slv_reg189(15 downto 0);
out_0_6 <= 		   slv_reg0(15 downto 0) * slv_reg134(15 downto 0)	 + slv_reg1(15 downto 0) * slv_reg142(15 downto 0)
				 + slv_reg2(15 downto 0) * slv_reg150(15 downto 0)	 + slv_reg3(15 downto 0) * slv_reg158(15 downto 0)
				 + slv_reg4(15 downto 0) * slv_reg166(15 downto 0)	 + slv_reg5(15 downto 0) * slv_reg174(15 downto 0)
				 + slv_reg6(15 downto 0) * slv_reg182(15 downto 0)	 + slv_reg7(15 downto 0) * slv_reg190(15 downto 0);
out_0_7 <= 		   slv_reg0(15 downto 0) * slv_reg135(15 downto 0)	 + slv_reg1(15 downto 0) * slv_reg143(15 downto 0)
				 + slv_reg2(15 downto 0) * slv_reg151(15 downto 0)	 + slv_reg3(15 downto 0) * slv_reg159(15 downto 0)
				 + slv_reg4(15 downto 0) * slv_reg167(15 downto 0)	 + slv_reg5(15 downto 0) * slv_reg175(15 downto 0)
				 + slv_reg6(15 downto 0) * slv_reg183(15 downto 0)	 + slv_reg7(15 downto 0) * slv_reg191(15 downto 0);
out_1_0 <= 		   slv_reg8(15 downto 0) * slv_reg128(15 downto 0)	 + slv_reg9(15 downto 0) * slv_reg136(15 downto 0)
				 + slv_reg10(15 downto 0) * slv_reg144(15 downto 0)	 + slv_reg11(15 downto 0) * slv_reg152(15 downto 0)
				 + slv_reg12(15 downto 0) * slv_reg160(15 downto 0)	 + slv_reg13(15 downto 0) * slv_reg168(15 downto 0)
				 + slv_reg14(15 downto 0) * slv_reg176(15 downto 0)	 + slv_reg15(15 downto 0) * slv_reg184(15 downto 0);
out_1_1 <= 		   slv_reg8(15 downto 0) * slv_reg129(15 downto 0)	 + slv_reg9(15 downto 0) * slv_reg137(15 downto 0)
				 + slv_reg10(15 downto 0) * slv_reg145(15 downto 0)	 + slv_reg11(15 downto 0) * slv_reg153(15 downto 0)
				 + slv_reg12(15 downto 0) * slv_reg161(15 downto 0)	 + slv_reg13(15 downto 0) * slv_reg169(15 downto 0)
				 + slv_reg14(15 downto 0) * slv_reg177(15 downto 0)	 + slv_reg15(15 downto 0) * slv_reg185(15 downto 0);
out_1_2 <= 		   slv_reg8(15 downto 0) * slv_reg130(15 downto 0)	 + slv_reg9(15 downto 0) * slv_reg138(15 downto 0)
				 + slv_reg10(15 downto 0) * slv_reg146(15 downto 0)	 + slv_reg11(15 downto 0) * slv_reg154(15 downto 0)
				 + slv_reg12(15 downto 0) * slv_reg162(15 downto 0)	 + slv_reg13(15 downto 0) * slv_reg170(15 downto 0)
				 + slv_reg14(15 downto 0) * slv_reg178(15 downto 0)	 + slv_reg15(15 downto 0) * slv_reg186(15 downto 0);
out_1_3 <= 		   slv_reg8(15 downto 0) * slv_reg131(15 downto 0)	 + slv_reg9(15 downto 0) * slv_reg139(15 downto 0)
				 + slv_reg10(15 downto 0) * slv_reg147(15 downto 0)	 + slv_reg11(15 downto 0) * slv_reg155(15 downto 0)
				 + slv_reg12(15 downto 0) * slv_reg163(15 downto 0)	 + slv_reg13(15 downto 0) * slv_reg171(15 downto 0)
				 + slv_reg14(15 downto 0) * slv_reg179(15 downto 0)	 + slv_reg15(15 downto 0) * slv_reg187(15 downto 0);
out_1_4 <= 		   slv_reg8(15 downto 0) * slv_reg132(15 downto 0)	 + slv_reg9(15 downto 0) * slv_reg140(15 downto 0)
				 + slv_reg10(15 downto 0) * slv_reg148(15 downto 0)	 + slv_reg11(15 downto 0) * slv_reg156(15 downto 0)
				 + slv_reg12(15 downto 0) * slv_reg164(15 downto 0)	 + slv_reg13(15 downto 0) * slv_reg172(15 downto 0)
				 + slv_reg14(15 downto 0) * slv_reg180(15 downto 0)	 + slv_reg15(15 downto 0) * slv_reg188(15 downto 0);
out_1_5 <= 		   slv_reg8(15 downto 0) * slv_reg133(15 downto 0)	 + slv_reg9(15 downto 0) * slv_reg141(15 downto 0)
				 + slv_reg10(15 downto 0) * slv_reg149(15 downto 0)	 + slv_reg11(15 downto 0) * slv_reg157(15 downto 0)
				 + slv_reg12(15 downto 0) * slv_reg165(15 downto 0)	 + slv_reg13(15 downto 0) * slv_reg173(15 downto 0)
				 + slv_reg14(15 downto 0) * slv_reg181(15 downto 0)	 + slv_reg15(15 downto 0) * slv_reg189(15 downto 0);
out_1_6 <= 		   slv_reg8(15 downto 0) * slv_reg134(15 downto 0)	 + slv_reg9(15 downto 0) * slv_reg142(15 downto 0)
				 + slv_reg10(15 downto 0) * slv_reg150(15 downto 0)	 + slv_reg11(15 downto 0) * slv_reg158(15 downto 0)
				 + slv_reg12(15 downto 0) * slv_reg166(15 downto 0)	 + slv_reg13(15 downto 0) * slv_reg174(15 downto 0)
				 + slv_reg14(15 downto 0) * slv_reg182(15 downto 0)	 + slv_reg15(15 downto 0) * slv_reg190(15 downto 0);
out_1_7 <= 		   slv_reg8(15 downto 0) * slv_reg135(15 downto 0)	 + slv_reg9(15 downto 0) * slv_reg143(15 downto 0)
				 + slv_reg10(15 downto 0) * slv_reg151(15 downto 0)	 + slv_reg11(15 downto 0) * slv_reg159(15 downto 0)
				 + slv_reg12(15 downto 0) * slv_reg167(15 downto 0)	 + slv_reg13(15 downto 0) * slv_reg175(15 downto 0)
				 + slv_reg14(15 downto 0) * slv_reg183(15 downto 0)	 + slv_reg15(15 downto 0) * slv_reg191(15 downto 0);
out_2_0 <= 		   slv_reg16(15 downto 0) * slv_reg128(15 downto 0)	 + slv_reg17(15 downto 0) * slv_reg136(15 downto 0)
				 + slv_reg18(15 downto 0) * slv_reg144(15 downto 0)	 + slv_reg19(15 downto 0) * slv_reg152(15 downto 0)
				 + slv_reg20(15 downto 0) * slv_reg160(15 downto 0)	 + slv_reg21(15 downto 0) * slv_reg168(15 downto 0)
				 + slv_reg22(15 downto 0) * slv_reg176(15 downto 0)	 + slv_reg23(15 downto 0) * slv_reg184(15 downto 0);
out_2_1 <= 		   slv_reg16(15 downto 0) * slv_reg129(15 downto 0)	 + slv_reg17(15 downto 0) * slv_reg137(15 downto 0)
				 + slv_reg18(15 downto 0) * slv_reg145(15 downto 0)	 + slv_reg19(15 downto 0) * slv_reg153(15 downto 0)
				 + slv_reg20(15 downto 0) * slv_reg161(15 downto 0)	 + slv_reg21(15 downto 0) * slv_reg169(15 downto 0)
				 + slv_reg22(15 downto 0) * slv_reg177(15 downto 0)	 + slv_reg23(15 downto 0) * slv_reg185(15 downto 0);
out_2_2 <= 		   slv_reg16(15 downto 0) * slv_reg130(15 downto 0)	 + slv_reg17(15 downto 0) * slv_reg138(15 downto 0)
				 + slv_reg18(15 downto 0) * slv_reg146(15 downto 0)	 + slv_reg19(15 downto 0) * slv_reg154(15 downto 0)
				 + slv_reg20(15 downto 0) * slv_reg162(15 downto 0)	 + slv_reg21(15 downto 0) * slv_reg170(15 downto 0)
				 + slv_reg22(15 downto 0) * slv_reg178(15 downto 0)	 + slv_reg23(15 downto 0) * slv_reg186(15 downto 0);
out_2_3 <= 		   slv_reg16(15 downto 0) * slv_reg131(15 downto 0)	 + slv_reg17(15 downto 0) * slv_reg139(15 downto 0)
				 + slv_reg18(15 downto 0) * slv_reg147(15 downto 0)	 + slv_reg19(15 downto 0) * slv_reg155(15 downto 0)
				 + slv_reg20(15 downto 0) * slv_reg163(15 downto 0)	 + slv_reg21(15 downto 0) * slv_reg171(15 downto 0)
				 + slv_reg22(15 downto 0) * slv_reg179(15 downto 0)	 + slv_reg23(15 downto 0) * slv_reg187(15 downto 0);
out_2_4 <= 		   slv_reg16(15 downto 0) * slv_reg132(15 downto 0)	 + slv_reg17(15 downto 0) * slv_reg140(15 downto 0)
				 + slv_reg18(15 downto 0) * slv_reg148(15 downto 0)	 + slv_reg19(15 downto 0) * slv_reg156(15 downto 0)
				 + slv_reg20(15 downto 0) * slv_reg164(15 downto 0)	 + slv_reg21(15 downto 0) * slv_reg172(15 downto 0)
				 + slv_reg22(15 downto 0) * slv_reg180(15 downto 0)	 + slv_reg23(15 downto 0) * slv_reg188(15 downto 0);
out_2_5 <= 		   slv_reg16(15 downto 0) * slv_reg133(15 downto 0)	 + slv_reg17(15 downto 0) * slv_reg141(15 downto 0)
				 + slv_reg18(15 downto 0) * slv_reg149(15 downto 0)	 + slv_reg19(15 downto 0) * slv_reg157(15 downto 0)
				 + slv_reg20(15 downto 0) * slv_reg165(15 downto 0)	 + slv_reg21(15 downto 0) * slv_reg173(15 downto 0)
				 + slv_reg22(15 downto 0) * slv_reg181(15 downto 0)	 + slv_reg23(15 downto 0) * slv_reg189(15 downto 0);
out_2_6 <= 		   slv_reg16(15 downto 0) * slv_reg134(15 downto 0)	 + slv_reg17(15 downto 0) * slv_reg142(15 downto 0)
				 + slv_reg18(15 downto 0) * slv_reg150(15 downto 0)	 + slv_reg19(15 downto 0) * slv_reg158(15 downto 0)
				 + slv_reg20(15 downto 0) * slv_reg166(15 downto 0)	 + slv_reg21(15 downto 0) * slv_reg174(15 downto 0)
				 + slv_reg22(15 downto 0) * slv_reg182(15 downto 0)	 + slv_reg23(15 downto 0) * slv_reg190(15 downto 0);
out_2_7 <= 		   slv_reg16(15 downto 0) * slv_reg135(15 downto 0)	 + slv_reg17(15 downto 0) * slv_reg143(15 downto 0)
				 + slv_reg18(15 downto 0) * slv_reg151(15 downto 0)	 + slv_reg19(15 downto 0) * slv_reg159(15 downto 0)
				 + slv_reg20(15 downto 0) * slv_reg167(15 downto 0)	 + slv_reg21(15 downto 0) * slv_reg175(15 downto 0)
				 + slv_reg22(15 downto 0) * slv_reg183(15 downto 0)	 + slv_reg23(15 downto 0) * slv_reg191(15 downto 0);
out_3_0 <= 		   slv_reg24(15 downto 0) * slv_reg128(15 downto 0)	 + slv_reg25(15 downto 0) * slv_reg136(15 downto 0)
				 + slv_reg26(15 downto 0) * slv_reg144(15 downto 0)	 + slv_reg27(15 downto 0) * slv_reg152(15 downto 0)
				 + slv_reg28(15 downto 0) * slv_reg160(15 downto 0)	 + slv_reg29(15 downto 0) * slv_reg168(15 downto 0)
				 + slv_reg30(15 downto 0) * slv_reg176(15 downto 0)	 + slv_reg31(15 downto 0) * slv_reg184(15 downto 0);
out_3_1 <= 		   slv_reg24(15 downto 0) * slv_reg129(15 downto 0)	 + slv_reg25(15 downto 0) * slv_reg137(15 downto 0)
				 + slv_reg26(15 downto 0) * slv_reg145(15 downto 0)	 + slv_reg27(15 downto 0) * slv_reg153(15 downto 0)
				 + slv_reg28(15 downto 0) * slv_reg161(15 downto 0)	 + slv_reg29(15 downto 0) * slv_reg169(15 downto 0)
				 + slv_reg30(15 downto 0) * slv_reg177(15 downto 0)	 + slv_reg31(15 downto 0) * slv_reg185(15 downto 0);
out_3_2 <= 		   slv_reg24(15 downto 0) * slv_reg130(15 downto 0)	 + slv_reg25(15 downto 0) * slv_reg138(15 downto 0)
				 + slv_reg26(15 downto 0) * slv_reg146(15 downto 0)	 + slv_reg27(15 downto 0) * slv_reg154(15 downto 0)
				 + slv_reg28(15 downto 0) * slv_reg162(15 downto 0)	 + slv_reg29(15 downto 0) * slv_reg170(15 downto 0)
				 + slv_reg30(15 downto 0) * slv_reg178(15 downto 0)	 + slv_reg31(15 downto 0) * slv_reg186(15 downto 0);
out_3_3 <= 		   slv_reg24(15 downto 0) * slv_reg131(15 downto 0)	 + slv_reg25(15 downto 0) * slv_reg139(15 downto 0)
				 + slv_reg26(15 downto 0) * slv_reg147(15 downto 0)	 + slv_reg27(15 downto 0) * slv_reg155(15 downto 0)
				 + slv_reg28(15 downto 0) * slv_reg163(15 downto 0)	 + slv_reg29(15 downto 0) * slv_reg171(15 downto 0)
				 + slv_reg30(15 downto 0) * slv_reg179(15 downto 0)	 + slv_reg31(15 downto 0) * slv_reg187(15 downto 0);
out_3_4 <= 		   slv_reg24(15 downto 0) * slv_reg132(15 downto 0)	 + slv_reg25(15 downto 0) * slv_reg140(15 downto 0)
				 + slv_reg26(15 downto 0) * slv_reg148(15 downto 0)	 + slv_reg27(15 downto 0) * slv_reg156(15 downto 0)
				 + slv_reg28(15 downto 0) * slv_reg164(15 downto 0)	 + slv_reg29(15 downto 0) * slv_reg172(15 downto 0)
				 + slv_reg30(15 downto 0) * slv_reg180(15 downto 0)	 + slv_reg31(15 downto 0) * slv_reg188(15 downto 0);
out_3_5 <= 		   slv_reg24(15 downto 0) * slv_reg133(15 downto 0)	 + slv_reg25(15 downto 0) * slv_reg141(15 downto 0)
				 + slv_reg26(15 downto 0) * slv_reg149(15 downto 0)	 + slv_reg27(15 downto 0) * slv_reg157(15 downto 0)
				 + slv_reg28(15 downto 0) * slv_reg165(15 downto 0)	 + slv_reg29(15 downto 0) * slv_reg173(15 downto 0)
				 + slv_reg30(15 downto 0) * slv_reg181(15 downto 0)	 + slv_reg31(15 downto 0) * slv_reg189(15 downto 0);
out_3_6 <= 		   slv_reg24(15 downto 0) * slv_reg134(15 downto 0)	 + slv_reg25(15 downto 0) * slv_reg142(15 downto 0)
				 + slv_reg26(15 downto 0) * slv_reg150(15 downto 0)	 + slv_reg27(15 downto 0) * slv_reg158(15 downto 0)
				 + slv_reg28(15 downto 0) * slv_reg166(15 downto 0)	 + slv_reg29(15 downto 0) * slv_reg174(15 downto 0)
				 + slv_reg30(15 downto 0) * slv_reg182(15 downto 0)	 + slv_reg31(15 downto 0) * slv_reg190(15 downto 0);
out_3_7 <= 		   slv_reg24(15 downto 0) * slv_reg135(15 downto 0)	 + slv_reg25(15 downto 0) * slv_reg143(15 downto 0)
				 + slv_reg26(15 downto 0) * slv_reg151(15 downto 0)	 + slv_reg27(15 downto 0) * slv_reg159(15 downto 0)
				 + slv_reg28(15 downto 0) * slv_reg167(15 downto 0)	 + slv_reg29(15 downto 0) * slv_reg175(15 downto 0)
				 + slv_reg30(15 downto 0) * slv_reg183(15 downto 0)	 + slv_reg31(15 downto 0) * slv_reg191(15 downto 0);
out_4_0 <= 		   slv_reg32(15 downto 0) * slv_reg128(15 downto 0)	 + slv_reg33(15 downto 0) * slv_reg136(15 downto 0)
				 + slv_reg34(15 downto 0) * slv_reg144(15 downto 0)	 + slv_reg35(15 downto 0) * slv_reg152(15 downto 0)
				 + slv_reg36(15 downto 0) * slv_reg160(15 downto 0)	 + slv_reg37(15 downto 0) * slv_reg168(15 downto 0)
				 + slv_reg38(15 downto 0) * slv_reg176(15 downto 0)	 + slv_reg39(15 downto 0) * slv_reg184(15 downto 0);
out_4_1 <= 		   slv_reg32(15 downto 0) * slv_reg129(15 downto 0)	 + slv_reg33(15 downto 0) * slv_reg137(15 downto 0)
				 + slv_reg34(15 downto 0) * slv_reg145(15 downto 0)	 + slv_reg35(15 downto 0) * slv_reg153(15 downto 0)
				 + slv_reg36(15 downto 0) * slv_reg161(15 downto 0)	 + slv_reg37(15 downto 0) * slv_reg169(15 downto 0)
				 + slv_reg38(15 downto 0) * slv_reg177(15 downto 0)	 + slv_reg39(15 downto 0) * slv_reg185(15 downto 0);
out_4_2 <= 		   slv_reg32(15 downto 0) * slv_reg130(15 downto 0)	 + slv_reg33(15 downto 0) * slv_reg138(15 downto 0)
				 + slv_reg34(15 downto 0) * slv_reg146(15 downto 0)	 + slv_reg35(15 downto 0) * slv_reg154(15 downto 0)
				 + slv_reg36(15 downto 0) * slv_reg162(15 downto 0)	 + slv_reg37(15 downto 0) * slv_reg170(15 downto 0)
				 + slv_reg38(15 downto 0) * slv_reg178(15 downto 0)	 + slv_reg39(15 downto 0) * slv_reg186(15 downto 0);
out_4_3 <= 		   slv_reg32(15 downto 0) * slv_reg131(15 downto 0)	 + slv_reg33(15 downto 0) * slv_reg139(15 downto 0)
				 + slv_reg34(15 downto 0) * slv_reg147(15 downto 0)	 + slv_reg35(15 downto 0) * slv_reg155(15 downto 0)
				 + slv_reg36(15 downto 0) * slv_reg163(15 downto 0)	 + slv_reg37(15 downto 0) * slv_reg171(15 downto 0)
				 + slv_reg38(15 downto 0) * slv_reg179(15 downto 0)	 + slv_reg39(15 downto 0) * slv_reg187(15 downto 0);
out_4_4 <= 		   slv_reg32(15 downto 0) * slv_reg132(15 downto 0)	 + slv_reg33(15 downto 0) * slv_reg140(15 downto 0)
				 + slv_reg34(15 downto 0) * slv_reg148(15 downto 0)	 + slv_reg35(15 downto 0) * slv_reg156(15 downto 0)
				 + slv_reg36(15 downto 0) * slv_reg164(15 downto 0)	 + slv_reg37(15 downto 0) * slv_reg172(15 downto 0)
				 + slv_reg38(15 downto 0) * slv_reg180(15 downto 0)	 + slv_reg39(15 downto 0) * slv_reg188(15 downto 0);
out_4_5 <= 		   slv_reg32(15 downto 0) * slv_reg133(15 downto 0)	 + slv_reg33(15 downto 0) * slv_reg141(15 downto 0)
				 + slv_reg34(15 downto 0) * slv_reg149(15 downto 0)	 + slv_reg35(15 downto 0) * slv_reg157(15 downto 0)
				 + slv_reg36(15 downto 0) * slv_reg165(15 downto 0)	 + slv_reg37(15 downto 0) * slv_reg173(15 downto 0)
				 + slv_reg38(15 downto 0) * slv_reg181(15 downto 0)	 + slv_reg39(15 downto 0) * slv_reg189(15 downto 0);
out_4_6 <= 		   slv_reg32(15 downto 0) * slv_reg134(15 downto 0)	 + slv_reg33(15 downto 0) * slv_reg142(15 downto 0)
				 + slv_reg34(15 downto 0) * slv_reg150(15 downto 0)	 + slv_reg35(15 downto 0) * slv_reg158(15 downto 0)
				 + slv_reg36(15 downto 0) * slv_reg166(15 downto 0)	 + slv_reg37(15 downto 0) * slv_reg174(15 downto 0)
				 + slv_reg38(15 downto 0) * slv_reg182(15 downto 0)	 + slv_reg39(15 downto 0) * slv_reg190(15 downto 0);
out_4_7 <= 		   slv_reg32(15 downto 0) * slv_reg135(15 downto 0)	 + slv_reg33(15 downto 0) * slv_reg143(15 downto 0)
				 + slv_reg34(15 downto 0) * slv_reg151(15 downto 0)	 + slv_reg35(15 downto 0) * slv_reg159(15 downto 0)
				 + slv_reg36(15 downto 0) * slv_reg167(15 downto 0)	 + slv_reg37(15 downto 0) * slv_reg175(15 downto 0)
				 + slv_reg38(15 downto 0) * slv_reg183(15 downto 0)	 + slv_reg39(15 downto 0) * slv_reg191(15 downto 0);
out_5_0 <= 		   slv_reg40(15 downto 0) * slv_reg128(15 downto 0)	 + slv_reg41(15 downto 0) * slv_reg136(15 downto 0)
				 + slv_reg42(15 downto 0) * slv_reg144(15 downto 0)	 + slv_reg43(15 downto 0) * slv_reg152(15 downto 0)
				 + slv_reg44(15 downto 0) * slv_reg160(15 downto 0)	 + slv_reg45(15 downto 0) * slv_reg168(15 downto 0)
				 + slv_reg46(15 downto 0) * slv_reg176(15 downto 0)	 + slv_reg47(15 downto 0) * slv_reg184(15 downto 0);
out_5_1 <= 		   slv_reg40(15 downto 0) * slv_reg129(15 downto 0)	 + slv_reg41(15 downto 0) * slv_reg137(15 downto 0)
				 + slv_reg42(15 downto 0) * slv_reg145(15 downto 0)	 + slv_reg43(15 downto 0) * slv_reg153(15 downto 0)
				 + slv_reg44(15 downto 0) * slv_reg161(15 downto 0)	 + slv_reg45(15 downto 0) * slv_reg169(15 downto 0)
				 + slv_reg46(15 downto 0) * slv_reg177(15 downto 0)	 + slv_reg47(15 downto 0) * slv_reg185(15 downto 0);
out_5_2 <= 		   slv_reg40(15 downto 0) * slv_reg130(15 downto 0)	 + slv_reg41(15 downto 0) * slv_reg138(15 downto 0)
				 + slv_reg42(15 downto 0) * slv_reg146(15 downto 0)	 + slv_reg43(15 downto 0) * slv_reg154(15 downto 0)
				 + slv_reg44(15 downto 0) * slv_reg162(15 downto 0)	 + slv_reg45(15 downto 0) * slv_reg170(15 downto 0)
				 + slv_reg46(15 downto 0) * slv_reg178(15 downto 0)	 + slv_reg47(15 downto 0) * slv_reg186(15 downto 0);
out_5_3 <= 		   slv_reg40(15 downto 0) * slv_reg131(15 downto 0)	 + slv_reg41(15 downto 0) * slv_reg139(15 downto 0)
				 + slv_reg42(15 downto 0) * slv_reg147(15 downto 0)	 + slv_reg43(15 downto 0) * slv_reg155(15 downto 0)
				 + slv_reg44(15 downto 0) * slv_reg163(15 downto 0)	 + slv_reg45(15 downto 0) * slv_reg171(15 downto 0)
				 + slv_reg46(15 downto 0) * slv_reg179(15 downto 0)	 + slv_reg47(15 downto 0) * slv_reg187(15 downto 0);
out_5_4 <= 		   slv_reg40(15 downto 0) * slv_reg132(15 downto 0)	 + slv_reg41(15 downto 0) * slv_reg140(15 downto 0)
				 + slv_reg42(15 downto 0) * slv_reg148(15 downto 0)	 + slv_reg43(15 downto 0) * slv_reg156(15 downto 0)
				 + slv_reg44(15 downto 0) * slv_reg164(15 downto 0)	 + slv_reg45(15 downto 0) * slv_reg172(15 downto 0)
				 + slv_reg46(15 downto 0) * slv_reg180(15 downto 0)	 + slv_reg47(15 downto 0) * slv_reg188(15 downto 0);
out_5_5 <= 		   slv_reg40(15 downto 0) * slv_reg133(15 downto 0)	 + slv_reg41(15 downto 0) * slv_reg141(15 downto 0)
				 + slv_reg42(15 downto 0) * slv_reg149(15 downto 0)	 + slv_reg43(15 downto 0) * slv_reg157(15 downto 0)
				 + slv_reg44(15 downto 0) * slv_reg165(15 downto 0)	 + slv_reg45(15 downto 0) * slv_reg173(15 downto 0)
				 + slv_reg46(15 downto 0) * slv_reg181(15 downto 0)	 + slv_reg47(15 downto 0) * slv_reg189(15 downto 0);
out_5_6 <= 		   slv_reg40(15 downto 0) * slv_reg134(15 downto 0)	 + slv_reg41(15 downto 0) * slv_reg142(15 downto 0)
				 + slv_reg42(15 downto 0) * slv_reg150(15 downto 0)	 + slv_reg43(15 downto 0) * slv_reg158(15 downto 0)
				 + slv_reg44(15 downto 0) * slv_reg166(15 downto 0)	 + slv_reg45(15 downto 0) * slv_reg174(15 downto 0)
				 + slv_reg46(15 downto 0) * slv_reg182(15 downto 0)	 + slv_reg47(15 downto 0) * slv_reg190(15 downto 0);
out_5_7 <= 		   slv_reg40(15 downto 0) * slv_reg135(15 downto 0)	 + slv_reg41(15 downto 0) * slv_reg143(15 downto 0)
				 + slv_reg42(15 downto 0) * slv_reg151(15 downto 0)	 + slv_reg43(15 downto 0) * slv_reg159(15 downto 0)
				 + slv_reg44(15 downto 0) * slv_reg167(15 downto 0)	 + slv_reg45(15 downto 0) * slv_reg175(15 downto 0)
				 + slv_reg46(15 downto 0) * slv_reg183(15 downto 0)	 + slv_reg47(15 downto 0) * slv_reg191(15 downto 0);
out_6_0 <= 		   slv_reg48(15 downto 0) * slv_reg128(15 downto 0)	 + slv_reg49(15 downto 0) * slv_reg136(15 downto 0)
				 + slv_reg50(15 downto 0) * slv_reg144(15 downto 0)	 + slv_reg51(15 downto 0) * slv_reg152(15 downto 0)
				 + slv_reg52(15 downto 0) * slv_reg160(15 downto 0)	 + slv_reg53(15 downto 0) * slv_reg168(15 downto 0)
				 + slv_reg54(15 downto 0) * slv_reg176(15 downto 0)	 + slv_reg55(15 downto 0) * slv_reg184(15 downto 0);
out_6_1 <= 		   slv_reg48(15 downto 0) * slv_reg129(15 downto 0)	 + slv_reg49(15 downto 0) * slv_reg137(15 downto 0)
				 + slv_reg50(15 downto 0) * slv_reg145(15 downto 0)	 + slv_reg51(15 downto 0) * slv_reg153(15 downto 0)
				 + slv_reg52(15 downto 0) * slv_reg161(15 downto 0)	 + slv_reg53(15 downto 0) * slv_reg169(15 downto 0)
				 + slv_reg54(15 downto 0) * slv_reg177(15 downto 0)	 + slv_reg55(15 downto 0) * slv_reg185(15 downto 0);
out_6_2 <= 		   slv_reg48(15 downto 0) * slv_reg130(15 downto 0)	 + slv_reg49(15 downto 0) * slv_reg138(15 downto 0)
				 + slv_reg50(15 downto 0) * slv_reg146(15 downto 0)	 + slv_reg51(15 downto 0) * slv_reg154(15 downto 0)
				 + slv_reg52(15 downto 0) * slv_reg162(15 downto 0)	 + slv_reg53(15 downto 0) * slv_reg170(15 downto 0)
				 + slv_reg54(15 downto 0) * slv_reg178(15 downto 0)	 + slv_reg55(15 downto 0) * slv_reg186(15 downto 0);
out_6_3 <= 		   slv_reg48(15 downto 0) * slv_reg131(15 downto 0)	 + slv_reg49(15 downto 0) * slv_reg139(15 downto 0)
				 + slv_reg50(15 downto 0) * slv_reg147(15 downto 0)	 + slv_reg51(15 downto 0) * slv_reg155(15 downto 0)
				 + slv_reg52(15 downto 0) * slv_reg163(15 downto 0)	 + slv_reg53(15 downto 0) * slv_reg171(15 downto 0)
				 + slv_reg54(15 downto 0) * slv_reg179(15 downto 0)	 + slv_reg55(15 downto 0) * slv_reg187(15 downto 0);
out_6_4 <= 		   slv_reg48(15 downto 0) * slv_reg132(15 downto 0)	 + slv_reg49(15 downto 0) * slv_reg140(15 downto 0)
				 + slv_reg50(15 downto 0) * slv_reg148(15 downto 0)	 + slv_reg51(15 downto 0) * slv_reg156(15 downto 0)
				 + slv_reg52(15 downto 0) * slv_reg164(15 downto 0)	 + slv_reg53(15 downto 0) * slv_reg172(15 downto 0)
				 + slv_reg54(15 downto 0) * slv_reg180(15 downto 0)	 + slv_reg55(15 downto 0) * slv_reg188(15 downto 0);
out_6_5 <= 		   slv_reg48(15 downto 0) * slv_reg133(15 downto 0)	 + slv_reg49(15 downto 0) * slv_reg141(15 downto 0)
				 + slv_reg50(15 downto 0) * slv_reg149(15 downto 0)	 + slv_reg51(15 downto 0) * slv_reg157(15 downto 0)
				 + slv_reg52(15 downto 0) * slv_reg165(15 downto 0)	 + slv_reg53(15 downto 0) * slv_reg173(15 downto 0)
				 + slv_reg54(15 downto 0) * slv_reg181(15 downto 0)	 + slv_reg55(15 downto 0) * slv_reg189(15 downto 0);
out_6_6 <= 		   slv_reg48(15 downto 0) * slv_reg134(15 downto 0)	 + slv_reg49(15 downto 0) * slv_reg142(15 downto 0)
				 + slv_reg50(15 downto 0) * slv_reg150(15 downto 0)	 + slv_reg51(15 downto 0) * slv_reg158(15 downto 0)
				 + slv_reg52(15 downto 0) * slv_reg166(15 downto 0)	 + slv_reg53(15 downto 0) * slv_reg174(15 downto 0)
				 + slv_reg54(15 downto 0) * slv_reg182(15 downto 0)	 + slv_reg55(15 downto 0) * slv_reg190(15 downto 0);
out_6_7 <= 		   slv_reg48(15 downto 0) * slv_reg135(15 downto 0)	 + slv_reg49(15 downto 0) * slv_reg143(15 downto 0)
				 + slv_reg50(15 downto 0) * slv_reg151(15 downto 0)	 + slv_reg51(15 downto 0) * slv_reg159(15 downto 0)
				 + slv_reg52(15 downto 0) * slv_reg167(15 downto 0)	 + slv_reg53(15 downto 0) * slv_reg175(15 downto 0)
				 + slv_reg54(15 downto 0) * slv_reg183(15 downto 0)	 + slv_reg55(15 downto 0) * slv_reg191(15 downto 0);
out_7_0 <= 		   slv_reg56(15 downto 0) * slv_reg128(15 downto 0)	 + slv_reg57(15 downto 0) * slv_reg136(15 downto 0)
				 + slv_reg58(15 downto 0) * slv_reg144(15 downto 0)	 + slv_reg59(15 downto 0) * slv_reg152(15 downto 0)
				 + slv_reg60(15 downto 0) * slv_reg160(15 downto 0)	 + slv_reg61(15 downto 0) * slv_reg168(15 downto 0)
				 + slv_reg62(15 downto 0) * slv_reg176(15 downto 0)	 + slv_reg63(15 downto 0) * slv_reg184(15 downto 0);
out_7_1 <= 		   slv_reg56(15 downto 0) * slv_reg129(15 downto 0)	 + slv_reg57(15 downto 0) * slv_reg137(15 downto 0)
				 + slv_reg58(15 downto 0) * slv_reg145(15 downto 0)	 + slv_reg59(15 downto 0) * slv_reg153(15 downto 0)
				 + slv_reg60(15 downto 0) * slv_reg161(15 downto 0)	 + slv_reg61(15 downto 0) * slv_reg169(15 downto 0)
				 + slv_reg62(15 downto 0) * slv_reg177(15 downto 0)	 + slv_reg63(15 downto 0) * slv_reg185(15 downto 0);
out_7_2 <= 		   slv_reg56(15 downto 0) * slv_reg130(15 downto 0)	 + slv_reg57(15 downto 0) * slv_reg138(15 downto 0)
				 + slv_reg58(15 downto 0) * slv_reg146(15 downto 0)	 + slv_reg59(15 downto 0) * slv_reg154(15 downto 0)
				 + slv_reg60(15 downto 0) * slv_reg162(15 downto 0)	 + slv_reg61(15 downto 0) * slv_reg170(15 downto 0)
				 + slv_reg62(15 downto 0) * slv_reg178(15 downto 0)	 + slv_reg63(15 downto 0) * slv_reg186(15 downto 0);
out_7_3 <= 		   slv_reg56(15 downto 0) * slv_reg131(15 downto 0)	 + slv_reg57(15 downto 0) * slv_reg139(15 downto 0)
				 + slv_reg58(15 downto 0) * slv_reg147(15 downto 0)	 + slv_reg59(15 downto 0) * slv_reg155(15 downto 0)
				 + slv_reg60(15 downto 0) * slv_reg163(15 downto 0)	 + slv_reg61(15 downto 0) * slv_reg171(15 downto 0)
				 + slv_reg62(15 downto 0) * slv_reg179(15 downto 0)	 + slv_reg63(15 downto 0) * slv_reg187(15 downto 0);
out_7_4 <= 		   slv_reg56(15 downto 0) * slv_reg132(15 downto 0)	 + slv_reg57(15 downto 0) * slv_reg140(15 downto 0)
				 + slv_reg58(15 downto 0) * slv_reg148(15 downto 0)	 + slv_reg59(15 downto 0) * slv_reg156(15 downto 0)
				 + slv_reg60(15 downto 0) * slv_reg164(15 downto 0)	 + slv_reg61(15 downto 0) * slv_reg172(15 downto 0)
				 + slv_reg62(15 downto 0) * slv_reg180(15 downto 0)	 + slv_reg63(15 downto 0) * slv_reg188(15 downto 0);
out_7_5 <= 		   slv_reg56(15 downto 0) * slv_reg133(15 downto 0)	 + slv_reg57(15 downto 0) * slv_reg141(15 downto 0)
				 + slv_reg58(15 downto 0) * slv_reg149(15 downto 0)	 + slv_reg59(15 downto 0) * slv_reg157(15 downto 0)
				 + slv_reg60(15 downto 0) * slv_reg165(15 downto 0)	 + slv_reg61(15 downto 0) * slv_reg173(15 downto 0)
				 + slv_reg62(15 downto 0) * slv_reg181(15 downto 0)	 + slv_reg63(15 downto 0) * slv_reg189(15 downto 0);
out_7_6 <= 		   slv_reg56(15 downto 0) * slv_reg134(15 downto 0)	 + slv_reg57(15 downto 0) * slv_reg142(15 downto 0)
				 + slv_reg58(15 downto 0) * slv_reg150(15 downto 0)	 + slv_reg59(15 downto 0) * slv_reg158(15 downto 0)
				 + slv_reg60(15 downto 0) * slv_reg166(15 downto 0)	 + slv_reg61(15 downto 0) * slv_reg174(15 downto 0)
				 + slv_reg62(15 downto 0) * slv_reg182(15 downto 0)	 + slv_reg63(15 downto 0) * slv_reg190(15 downto 0);
out_7_7 <= 		   slv_reg56(15 downto 0) * slv_reg135(15 downto 0)	 + slv_reg57(15 downto 0) * slv_reg143(15 downto 0)
				 + slv_reg58(15 downto 0) * slv_reg151(15 downto 0)	 + slv_reg59(15 downto 0) * slv_reg159(15 downto 0)
				 + slv_reg60(15 downto 0) * slv_reg167(15 downto 0)	 + slv_reg61(15 downto 0) * slv_reg175(15 downto 0)
				 + slv_reg62(15 downto 0) * slv_reg183(15 downto 0)	 + slv_reg63(15 downto 0) * slv_reg191(15 downto 0);


--  = # = # = # = # = # = # = # = # = # = # = # = # = # = # = # = # = # = # = # = # = # = # = # = # = # = # = # = #
--  = # = # = # = # = # = # = # = # = # = # = # = # = # = # = # = # = # = # = # = # = # = # = # = # = # = # = # = #


--                          R E G I S T E R    A C C E S S



process (slv_reg0, slv_reg1, slv_reg2, slv_reg3, slv_reg4, slv_reg5, slv_reg6, slv_reg7, slv_reg8, slv_reg9, slv_reg10, slv_reg11, slv_reg12, slv_reg13, slv_reg14, slv_reg15, slv_reg16, slv_reg17, slv_reg18, slv_reg19, slv_reg20, slv_reg21, slv_reg22, slv_reg23, slv_reg24, slv_reg25, slv_reg26, slv_reg27, slv_reg28, slv_reg29, slv_reg30, slv_reg31, slv_reg32, slv_reg33, slv_reg34, slv_reg35, slv_reg36, slv_reg37, slv_reg38, slv_reg39, slv_reg40, slv_reg41, slv_reg42, slv_reg43, slv_reg44, slv_reg45, slv_reg46, slv_reg47, slv_reg48, slv_reg49, slv_reg50, slv_reg51, slv_reg52, slv_reg53, slv_reg54, slv_reg55, slv_reg56, slv_reg57, slv_reg58, slv_reg59, slv_reg60, slv_reg61, slv_reg62, slv_reg63, slv_reg64, slv_reg65, slv_reg66, slv_reg67, slv_reg68, slv_reg69, slv_reg70, slv_reg71, slv_reg72, slv_reg73, slv_reg74, slv_reg75, slv_reg76, slv_reg77, slv_reg78, slv_reg79, slv_reg80, slv_reg81, slv_reg82, slv_reg83, slv_reg84, slv_reg85, slv_reg86, slv_reg87, slv_reg88, slv_reg89, slv_reg90, slv_reg91, slv_reg92, slv_reg93, slv_reg94, slv_reg95, slv_reg96, slv_reg97, slv_reg98, slv_reg99, slv_reg100, slv_reg101, slv_reg102, slv_reg103, slv_reg104, slv_reg105, slv_reg106, slv_reg107, slv_reg108, slv_reg109, slv_reg110, slv_reg111, slv_reg112, slv_reg113, slv_reg114, slv_reg115, slv_reg116, slv_reg117, slv_reg118, slv_reg119, slv_reg120, slv_reg121, slv_reg122, slv_reg123, slv_reg124, slv_reg125, slv_reg126, slv_reg127, slv_reg128, slv_reg129, slv_reg130, slv_reg131, slv_reg132, slv_reg133, slv_reg134, slv_reg135, slv_reg136, slv_reg137, slv_reg138, slv_reg139, slv_reg140, slv_reg141, slv_reg142, slv_reg143, slv_reg144, slv_reg145, slv_reg146, slv_reg147, slv_reg148, slv_reg149, slv_reg150, slv_reg151, slv_reg152, slv_reg153, slv_reg154, slv_reg155, slv_reg156, slv_reg157, slv_reg158, slv_reg159, slv_reg160, slv_reg161, slv_reg162, slv_reg163, slv_reg164, slv_reg165, slv_reg166, slv_reg167, slv_reg168, slv_reg169, slv_reg170, slv_reg171, slv_reg172, slv_reg173, slv_reg174, slv_reg175, slv_reg176, slv_reg177, slv_reg178, slv_reg179, slv_reg180, slv_reg181, slv_reg182, slv_reg183, slv_reg184, slv_reg185, slv_reg186, slv_reg187, slv_reg188, slv_reg189, slv_reg190, slv_reg191, slv_reg192, slv_reg193, slv_reg194, slv_reg195, slv_reg196, slv_reg197, slv_reg198, slv_reg199, slv_reg200, slv_reg201, slv_reg202, slv_reg203, slv_reg204, slv_reg205, slv_reg206, slv_reg207, slv_reg208, slv_reg209, slv_reg210, slv_reg211, slv_reg212, slv_reg213, slv_reg214, slv_reg215, slv_reg216, slv_reg217, slv_reg218, slv_reg219, slv_reg220, slv_reg221, slv_reg222, slv_reg223, slv_reg224, slv_reg225, slv_reg226, slv_reg227, slv_reg228, slv_reg229, slv_reg230, slv_reg231, slv_reg232, slv_reg233, slv_reg234, slv_reg235, slv_reg236, slv_reg237, slv_reg238, slv_reg239, slv_reg240, slv_reg241, slv_reg242, slv_reg243, slv_reg244, slv_reg245, slv_reg246, slv_reg247, slv_reg248, slv_reg249, slv_reg250, slv_reg251, slv_reg252, slv_reg253, slv_reg254, slv_reg255, slv_reg256, slv_reg257, slv_reg258, slv_reg259, slv_reg260, slv_reg261, slv_reg262, slv_reg263, slv_reg264, slv_reg265, slv_reg266, slv_reg267, slv_reg268, slv_reg269, slv_reg270, slv_reg271, slv_reg272, slv_reg273, slv_reg274, slv_reg275, slv_reg276, slv_reg277, slv_reg278, slv_reg279, slv_reg280, slv_reg281, slv_reg282, slv_reg283, slv_reg284, slv_reg285, slv_reg286, slv_reg287, slv_reg288, slv_reg289, slv_reg290, slv_reg291, slv_reg292, slv_reg293, slv_reg294, slv_reg295, slv_reg296, slv_reg297, slv_reg298, slv_reg299, slv_reg300, slv_reg301, slv_reg302, slv_reg303, slv_reg304, slv_reg305, slv_reg306, slv_reg307, slv_reg308, slv_reg309, slv_reg310, slv_reg311, slv_reg312, slv_reg313, slv_reg314, slv_reg315, slv_reg316, slv_reg317, slv_reg318, slv_reg319, slv_reg320, slv_reg321, slv_reg322, slv_reg323, slv_reg324, slv_reg325, slv_reg326, slv_reg327, slv_reg328, slv_reg329, slv_reg330, slv_reg331, slv_reg332, slv_reg333, slv_reg334, slv_reg335, slv_reg336, slv_reg337, slv_reg338, slv_reg339, slv_reg340, slv_reg341, slv_reg342, slv_reg343, slv_reg344, slv_reg345, slv_reg346, slv_reg347, slv_reg348, slv_reg349, slv_reg350, slv_reg351, slv_reg352, slv_reg353, slv_reg354, slv_reg355, slv_reg356, slv_reg357, slv_reg358, slv_reg359, slv_reg360, slv_reg361, slv_reg362, slv_reg363, slv_reg364, slv_reg365, slv_reg366, slv_reg367, slv_reg368, slv_reg369, slv_reg370, slv_reg371, slv_reg372, slv_reg373, slv_reg374, slv_reg375, slv_reg376, slv_reg377, slv_reg378, slv_reg379, slv_reg380, slv_reg381, slv_reg382, slv_reg383, slv_reg384, slv_reg385, slv_reg386, slv_reg387, slv_reg388, slv_reg389, slv_reg390, slv_reg391, slv_reg392, slv_reg393, slv_reg394, slv_reg395, slv_reg396, slv_reg397, slv_reg398, slv_reg399, slv_reg400, slv_reg401, slv_reg402, slv_reg403, slv_reg404, slv_reg405, slv_reg406, slv_reg407, slv_reg408, slv_reg409, slv_reg410, slv_reg411, slv_reg412, slv_reg413, slv_reg414, slv_reg415, slv_reg416, slv_reg417, slv_reg418, slv_reg419, slv_reg420, slv_reg421, slv_reg422, slv_reg423, slv_reg424, slv_reg425, slv_reg426, slv_reg427, slv_reg428, slv_reg429, slv_reg430, slv_reg431, slv_reg432, slv_reg433, slv_reg434, slv_reg435, slv_reg436, slv_reg437, slv_reg438, slv_reg439, slv_reg440, slv_reg441, slv_reg442, slv_reg443, slv_reg444, slv_reg445, slv_reg446, slv_reg447, slv_reg448, slv_reg449, slv_reg450, slv_reg451, slv_reg452, slv_reg453, slv_reg454, slv_reg455, slv_reg456, slv_reg457, slv_reg458, slv_reg459, slv_reg460, slv_reg461, slv_reg462, slv_reg463, slv_reg464, slv_reg465, slv_reg466, slv_reg467, slv_reg468, slv_reg469, slv_reg470, slv_reg471, slv_reg472, slv_reg473, slv_reg474, slv_reg475, slv_reg476, slv_reg477, slv_reg478, slv_reg479, slv_reg480, slv_reg481, slv_reg482, slv_reg483, slv_reg484, slv_reg485, slv_reg486, slv_reg487, slv_reg488, slv_reg489, slv_reg490, slv_reg491, slv_reg492, slv_reg493, slv_reg494, slv_reg495, slv_reg496, slv_reg497, slv_reg498, slv_reg499, slv_reg500, slv_reg501, slv_reg502, slv_reg503, slv_reg504, slv_reg505, slv_reg506, slv_reg507, slv_reg508, slv_reg509, slv_reg510, slv_reg511, axi_araddr, S_AXI_ARESETN, slv_reg_rden)
variable loc_addr :std_logic_vector(OPT_MEM_ADDR_BITS downto 0);
begin
loc_addr := axi_araddr(ADDR_LSB + OPT_MEM_ADDR_BITS downto ADDR_LSB);
    case loc_addr is
    
--  = # = # = # = # = # = # = # = # = # = # = # = # = # = # = # = # = # = # = # = # = # = # = # = # = # = # = # = #


    --  Control Signal   
 

    --  A Input
    
    when b"000000000" =>reg_data_out <= slv_reg0;      when b"000000001" =>reg_data_out <= slv_reg1;	
    when b"000000010" =>reg_data_out <= slv_reg2;      when b"000000011" =>reg_data_out <= slv_reg3;    
    when b"000000100" =>reg_data_out <= slv_reg4;      when b"000000101" =>reg_data_out <= slv_reg5;    
    when b"000000110" =>reg_data_out <= slv_reg6;      when b"000000111" =>reg_data_out <= slv_reg7;    
    when b"000001000" =>reg_data_out <= slv_reg8;      when b"000001001" =>reg_data_out <= slv_reg9;    
    when b"000001010" =>reg_data_out <= slv_reg10;     when b"000001011" =>reg_data_out <= slv_reg11;    
    when b"000001100" =>reg_data_out <= slv_reg12;     when b"000001101" =>reg_data_out <= slv_reg13;    
    when b"000001110" =>reg_data_out <= slv_reg14;     when b"000001111" =>reg_data_out <= slv_reg15;    
    when b"000010000" =>reg_data_out <= slv_reg16;     when b"000010001" =>reg_data_out <= slv_reg17;    
    when b"000010010" =>reg_data_out <= slv_reg18;     when b"000010011" =>reg_data_out <= slv_reg19;    
    when b"000010100" =>reg_data_out <= slv_reg20;     when b"000010101" =>reg_data_out <= slv_reg21;    
    when b"000010110" =>reg_data_out <= slv_reg22;     when b"000010111" =>reg_data_out <= slv_reg23;    
    when b"000011000" =>reg_data_out <= slv_reg24;     when b"000011001" =>reg_data_out <= slv_reg25;    
    when b"000011010" =>reg_data_out <= slv_reg26;     when b"000011011" =>reg_data_out <= slv_reg27;    
    when b"000011100" =>reg_data_out <= slv_reg28;     when b"000011101" =>reg_data_out <= slv_reg29;    
    when b"000011110" =>reg_data_out <= slv_reg30;     when b"000011111" =>reg_data_out <= slv_reg31;    
    when b"000100000" =>reg_data_out <= slv_reg32;     when b"000100001" =>reg_data_out <= slv_reg33;    
    when b"000100010" =>reg_data_out <= slv_reg34;     when b"000100011" =>reg_data_out <= slv_reg35;    
    when b"000100100" =>reg_data_out <= slv_reg36;     when b"000100101" =>reg_data_out <= slv_reg37;    
    when b"000100110" =>reg_data_out <= slv_reg38;     when b"000100111" =>reg_data_out <= slv_reg39;    
    when b"000101000" =>reg_data_out <= slv_reg40;     when b"000101001" =>reg_data_out <= slv_reg41;    
    when b"000101010" =>reg_data_out <= slv_reg42;     when b"000101011" =>reg_data_out <= slv_reg43;    
    when b"000101100" =>reg_data_out <= slv_reg44;     when b"000101101" =>reg_data_out <= slv_reg45;    
    when b"000101110" =>reg_data_out <= slv_reg46;     when b"000101111" =>reg_data_out <= slv_reg47;    
    when b"000110000" =>reg_data_out <= slv_reg48;     when b"000110001" =>reg_data_out <= slv_reg49;    
    when b"000110010" =>reg_data_out <= slv_reg50;     when b"000110011" =>reg_data_out <= slv_reg51;    
    when b"000110100" =>reg_data_out <= slv_reg52;     when b"000110101" =>reg_data_out <= slv_reg53;    
    when b"000110110" =>reg_data_out <= slv_reg54;     when b"000110111" =>reg_data_out <= slv_reg55;    
    when b"000111000" =>reg_data_out <= slv_reg56;     when b"000111001" =>reg_data_out <= slv_reg57;    
    when b"000111010" =>reg_data_out <= slv_reg58;     when b"000111011" =>reg_data_out <= slv_reg59;    
    when b"000111100" =>reg_data_out <= slv_reg60;     when b"000111101" =>reg_data_out <= slv_reg61;    
    when b"000111110" =>reg_data_out <= slv_reg62;     when b"000111111" =>reg_data_out <= slv_reg63;    
    when b"001000000" =>reg_data_out <= slv_reg64;     when b"001000001" =>reg_data_out <= slv_reg65;    
    when b"001000010" =>reg_data_out <= slv_reg66;     when b"001000011" =>reg_data_out <= slv_reg67;    
    when b"001000100" =>reg_data_out <= slv_reg68;     when b"001000101" =>reg_data_out <= slv_reg69;    
    when b"001000110" =>reg_data_out <= slv_reg70;     when b"001000111" =>reg_data_out <= slv_reg71;    
    when b"001001000" =>reg_data_out <= slv_reg72;     when b"001001001" =>reg_data_out <= slv_reg73;    
    when b"001001010" =>reg_data_out <= slv_reg74;     when b"001001011" =>reg_data_out <= slv_reg75;    
    when b"001001100" =>reg_data_out <= slv_reg76;     when b"001001101" =>reg_data_out <= slv_reg77;    
    when b"001001110" =>reg_data_out <= slv_reg78;     when b"001001111" =>reg_data_out <= slv_reg79;    
    when b"001010000" =>reg_data_out <= slv_reg80;     when b"001010001" =>reg_data_out <= slv_reg81;    
    when b"001010010" =>reg_data_out <= slv_reg82;     when b"001010011" =>reg_data_out <= slv_reg83;    
    when b"001010100" =>reg_data_out <= slv_reg84;     when b"001010101" =>reg_data_out <= slv_reg85;    
    when b"001010110" =>reg_data_out <= slv_reg86;     when b"001010111" =>reg_data_out <= slv_reg87;    
    when b"001011000" =>reg_data_out <= slv_reg88;     when b"001011001" =>reg_data_out <= slv_reg89;    
    when b"001011010" =>reg_data_out <= slv_reg90;     when b"001011011" =>reg_data_out <= slv_reg91;    
    when b"001011100" =>reg_data_out <= slv_reg92;     when b"001011101" =>reg_data_out <= slv_reg93;    
    when b"001011110" =>reg_data_out <= slv_reg94;     when b"001011111" =>reg_data_out <= slv_reg95;    
    when b"001100000" =>reg_data_out <= slv_reg96;     when b"001100001" =>reg_data_out <= slv_reg97;
    when b"001100010" =>reg_data_out <= slv_reg98;     when b"001100011" =>reg_data_out <= slv_reg99;    
    when b"001100100" =>reg_data_out <= slv_reg100;    when b"001100101" =>reg_data_out <= slv_reg101;    
    when b"001100110" =>reg_data_out <= slv_reg102;    when b"001100111" =>reg_data_out <= slv_reg103;    
    when b"001101000" =>reg_data_out <= slv_reg104;    when b"001101001" =>reg_data_out <= slv_reg105;    
    when b"001101010" =>reg_data_out <= slv_reg106;    when b"001101011" =>reg_data_out <= slv_reg107;    
    when b"001101100" =>reg_data_out <= slv_reg108;    when b"001101101" =>reg_data_out <= slv_reg109;    
    when b"001101110" =>reg_data_out <= slv_reg110;    when b"001101111" =>reg_data_out <= slv_reg111;    
    when b"001110000" =>reg_data_out <= slv_reg112;    when b"001110001" =>reg_data_out <= slv_reg113;    
    when b"001110010" =>reg_data_out <= slv_reg114;    when b"001110011" =>reg_data_out <= slv_reg115;    
    when b"001110100" =>reg_data_out <= slv_reg116;    when b"001110101" =>reg_data_out <= slv_reg117;    
    when b"001110110" =>reg_data_out <= slv_reg118;    when b"001110111" =>reg_data_out <= slv_reg119;    
    when b"001111000" =>reg_data_out <= slv_reg120;    when b"001111001" =>reg_data_out <= slv_reg121;    
    when b"001111010" =>reg_data_out <= slv_reg122;    when b"001111011" =>reg_data_out <= slv_reg123;    
    when b"001111100" =>reg_data_out <= slv_reg124;    when b"001111101" =>reg_data_out <= slv_reg125;    
    when b"001111110" =>reg_data_out <= slv_reg126;    when b"001111111" =>reg_data_out <= slv_reg127;
    
--  = # = # = # = # = # = # = # = # = # = # = # = # = # = # = # = # = # = # = # = # = # = # = # = # = # = # = # = #

--      B Input 
            
    when b"010000000" =>reg_data_out <= slv_reg128;    when b"010000001" =>reg_data_out <= slv_reg129;    
    when b"010000010" =>reg_data_out <= slv_reg130;    when b"010000011" =>reg_data_out <= slv_reg131;    
    when b"010000100" =>reg_data_out <= slv_reg132;    when b"010000101" =>reg_data_out <= slv_reg133;    
    when b"010000110" =>reg_data_out <= slv_reg134;    when b"010000111" =>reg_data_out <= slv_reg135;    
    when b"010001000" =>reg_data_out <= slv_reg136;    when b"010001001" =>reg_data_out <= slv_reg137;    
    when b"010001010" =>reg_data_out <= slv_reg138;    when b"010001011" =>reg_data_out <= slv_reg139;    
    when b"010001100" =>reg_data_out <= slv_reg140;    when b"010001101" =>reg_data_out <= slv_reg141;    
    when b"010001110" =>reg_data_out <= slv_reg142;    when b"010001111" =>reg_data_out <= slv_reg143;    
    when b"010010000" =>reg_data_out <= slv_reg144;    when b"010010001" =>reg_data_out <= slv_reg145;    
    when b"010010010" =>reg_data_out <= slv_reg146;    when b"010010011" =>reg_data_out <= slv_reg147;    
    when b"010010100" =>reg_data_out <= slv_reg148;    when b"010010101" =>reg_data_out <= slv_reg149;    
    when b"010010110" =>reg_data_out <= slv_reg150;    when b"010010111" =>reg_data_out <= slv_reg151;    
    when b"010011000" =>reg_data_out <= slv_reg152;    when b"010011001" =>reg_data_out <= slv_reg153;    
    when b"010011010" =>reg_data_out <= slv_reg154;    when b"010011011" =>reg_data_out <= slv_reg155;    
    when b"010011100" =>reg_data_out <= slv_reg156;    when b"010011101" =>reg_data_out <= slv_reg157;    
    when b"010011110" =>reg_data_out <= slv_reg158;    when b"010011111" =>reg_data_out <= slv_reg159;    
    when b"010100000" =>reg_data_out <= slv_reg160;    when b"010100001" =>reg_data_out <= slv_reg161;    
    when b"010100010" =>reg_data_out <= slv_reg162;    when b"010100011" =>reg_data_out <= slv_reg163;    
    when b"010100100" =>reg_data_out <= slv_reg164;    when b"010100101" =>reg_data_out <= slv_reg165;    
    when b"010100110" =>reg_data_out <= slv_reg166;    when b"010100111" =>reg_data_out <= slv_reg167;    
    when b"010101000" =>reg_data_out <= slv_reg168;    when b"010101001" =>reg_data_out <= slv_reg169;    
    when b"010101010" =>reg_data_out <= slv_reg170;    when b"010101011" =>reg_data_out <= slv_reg171;    
    when b"010101100" =>reg_data_out <= slv_reg172;    when b"010101101" =>reg_data_out <= slv_reg173;    
    when b"010101110" =>reg_data_out <= slv_reg174;    when b"010101111" =>reg_data_out <= slv_reg175;    
    when b"010110000" =>reg_data_out <= slv_reg176;    when b"010110001" =>reg_data_out <= slv_reg177;    
    when b"010110010" =>reg_data_out <= slv_reg178;    when b"010110011" =>reg_data_out <= slv_reg179;    
    when b"010110100" =>reg_data_out <= slv_reg180;    when b"010110101" =>reg_data_out <= slv_reg181;    
    when b"010110110" =>reg_data_out <= slv_reg182;    when b"010110111" =>reg_data_out <= slv_reg183;    
    when b"010111000" =>reg_data_out <= slv_reg184;    when b"010111001" =>reg_data_out <= slv_reg185;    
    when b"010111010" =>reg_data_out <= slv_reg186;    when b"010111011" =>reg_data_out <= slv_reg187;    
    when b"010111100" =>reg_data_out <= slv_reg188;    when b"010111101" =>reg_data_out <= slv_reg189;    
    when b"010111110" =>reg_data_out <= slv_reg190;    when b"010111111" =>reg_data_out <= slv_reg191;    
    when b"011000000" =>reg_data_out <= slv_reg192;    when b"011000001" =>reg_data_out <= slv_reg193;    
    when b"011000010" =>reg_data_out <= slv_reg194;    when b"011000011" =>reg_data_out <= slv_reg195;    
    when b"011000100" =>reg_data_out <= slv_reg196;    when b"011000101" =>reg_data_out <= slv_reg197;    
    when b"011000110" =>reg_data_out <= slv_reg198;    when b"011000111" =>reg_data_out <= slv_reg199;    
    when b"011001000" =>reg_data_out <= slv_reg200;    when b"011001001" =>reg_data_out <= slv_reg201;    
    when b"011001010" =>reg_data_out <= slv_reg202;    when b"011001011" =>reg_data_out <= slv_reg203;    
    when b"011001100" =>reg_data_out <= slv_reg204;    when b"011001101" =>reg_data_out <= slv_reg205;    
    when b"011001110" =>reg_data_out <= slv_reg206;    when b"011001111" =>reg_data_out <= slv_reg207;    
    when b"011010000" =>reg_data_out <= slv_reg208;    when b"011010001" =>reg_data_out <= slv_reg209;    
    when b"011010010" =>reg_data_out <= slv_reg210;    when b"011010011" =>reg_data_out <= slv_reg211;    
    when b"011010100" =>reg_data_out <= slv_reg212;    when b"011010101" =>reg_data_out <= slv_reg213;    
    when b"011010110" =>reg_data_out <= slv_reg214;    when b"011010111" =>reg_data_out <= slv_reg215;    
    when b"011011000" =>reg_data_out <= slv_reg216;    when b"011011001" =>reg_data_out <= slv_reg217;    
    when b"011011010" =>reg_data_out <= slv_reg218;    when b"011011011" =>reg_data_out <= slv_reg219;    
    when b"011011100" =>reg_data_out <= slv_reg220;    when b"011011101" =>reg_data_out <= slv_reg221;    
    when b"011011110" =>reg_data_out <= slv_reg222;    when b"011011111" =>reg_data_out <= slv_reg223;    
    when b"011100000" =>reg_data_out <= slv_reg224;    when b"011100001" =>reg_data_out <= slv_reg225;        
    when b"011100010" =>reg_data_out <= slv_reg226;    when b"011100011" =>reg_data_out <= slv_reg227;    
    when b"011100100" =>reg_data_out <= slv_reg228;    when b"011100101" =>reg_data_out <= slv_reg229;    
    when b"011100110" =>reg_data_out <= slv_reg230;    when b"011100111" =>reg_data_out <= slv_reg231;    
    when b"011101000" =>reg_data_out <= slv_reg232;    when b"011101001" =>reg_data_out <= slv_reg233;    
    when b"011101010" =>reg_data_out <= slv_reg234;    when b"011101011" =>reg_data_out <= slv_reg235;    
    when b"011101100" =>reg_data_out <= slv_reg236;    when b"011101101" =>reg_data_out <= slv_reg237;    
    when b"011101110" =>reg_data_out <= slv_reg238;    when b"011101111" =>reg_data_out <= slv_reg239;    
    when b"011110000" =>reg_data_out <= slv_reg240;    when b"011110001" =>reg_data_out <= slv_reg241;    
    when b"011110010" =>reg_data_out <= slv_reg242;    when b"011110011" =>reg_data_out <= slv_reg243;    
    when b"011110100" =>reg_data_out <= slv_reg244;    when b"011110101" =>reg_data_out <= slv_reg245;    
    when b"011110110" =>reg_data_out <= slv_reg246;    when b"011110111" =>reg_data_out <= slv_reg247;    
    when b"011111000" =>reg_data_out <= slv_reg248;    when b"011111001" =>reg_data_out <= slv_reg249;    
    when b"011111010" =>reg_data_out <= slv_reg250;    when b"011111011" =>reg_data_out <= slv_reg251;    
    when b"011111100" =>reg_data_out <= slv_reg252;    when b"011111101" =>reg_data_out <= slv_reg253;    
    when b"011111110" =>reg_data_out <= slv_reg254;    when b"011111111" =>reg_data_out <= slv_reg255;
    
--  = # = # = # = # = # = # = # = # = # = # = # = # = # = # = # = # = # = # = # = # = # = # = # = # = # = # = # = #

    --  C Output 
      
           
    when b"100000000" =>reg_data_out <= out_0_0;        when b"100000001"=>reg_data_out <= out_0_1;
    when b"100000010" =>reg_data_out <= out_0_2;        when b"100000011"=>reg_data_out <= out_0_3;
    when b"100000100" =>reg_data_out <= out_0_4;        when b"100000101"=>reg_data_out <= out_0_5;
    when b"100000110" =>reg_data_out <= out_0_6;        when b"100000111"=>reg_data_out <= out_0_7;
    when b"100001000" =>reg_data_out <= out_1_0;        when b"100001001"=>reg_data_out <= out_1_1;
    when b"100001010" =>reg_data_out <= out_1_2;        when b"100001011"=>reg_data_out <= out_1_3;
    when b"100001100" =>reg_data_out <= out_1_4;        when b"100001101"=>reg_data_out <= out_1_5;
    when b"100001110" =>reg_data_out <= out_1_6;        when b"100001111"=>reg_data_out <= out_1_7;
    when b"100010000" =>reg_data_out <= out_2_0;        when b"100010001"=>reg_data_out <= out_2_1;
    when b"100010010" =>reg_data_out <= out_2_2;        when b"100010011"=>reg_data_out <= out_2_3;
    when b"100010100" =>reg_data_out <= out_2_4;        when b"100010101"=>reg_data_out <= out_2_5;
    when b"100010110" =>reg_data_out <= out_2_6;        when b"100010111"=>reg_data_out <= out_2_7;
    when b"100011000" =>reg_data_out <= out_3_0;        when b"100011001"=>reg_data_out <= out_3_1;
    when b"100011010" =>reg_data_out <= out_3_2;        when b"100011011"=>reg_data_out <= out_3_3;
    when b"100011100" =>reg_data_out <= out_3_4;        when b"100011101"=>reg_data_out <= out_3_5;
    when b"100011110" =>reg_data_out <= out_3_6;        when b"100011111"=>reg_data_out <= out_3_7;
    when b"100100000" =>reg_data_out <= out_4_0;        when b"100100001"=>reg_data_out <= out_4_1;
    when b"100100010" =>reg_data_out <= out_4_2;        when b"100100011"=>reg_data_out <= out_4_3;
    when b"100100100" =>reg_data_out <= out_4_4;        when b"100100101"=>reg_data_out <= out_4_5;
    when b"100100110" =>reg_data_out <= out_4_6;        when b"100100111"=>reg_data_out <= out_4_7;
    when b"100101000" =>reg_data_out <= out_5_0;        when b"100101001"=>reg_data_out <= out_5_1;
    when b"100101010" =>reg_data_out <= out_5_2;        when b"100101011"=>reg_data_out <= out_5_3;
    when b"100101100" =>reg_data_out <= out_5_4;        when b"100101101"=>reg_data_out <= out_5_5;
    when b"100101110" =>reg_data_out <= out_5_6;        when b"100101111"=>reg_data_out <= out_5_7;
    when b"100110000" =>reg_data_out <= out_6_0;        when b"100110001"=>reg_data_out <= out_6_1;
    when b"100110010" =>reg_data_out <= out_6_2;        when b"100110011"=>reg_data_out <= out_6_3;
    when b"100110100" =>reg_data_out <= out_6_4;        when b"100110101"=>reg_data_out <= out_6_5;
    when b"100110110" =>reg_data_out <= out_6_6;        when b"100110111"=>reg_data_out <= out_6_7;
    when b"100111000" =>reg_data_out <= out_7_0;        when b"100111001"=>reg_data_out <= out_7_1;
    when b"100111010" =>reg_data_out <= out_7_2;        when b"100111011"=>reg_data_out <= out_7_3;
    when b"100111100" =>reg_data_out <= out_7_4;        when b"100111101"=>reg_data_out <= out_7_5;
    when b"100111110" =>reg_data_out <= out_7_6;        when b"100111111"=>reg_data_out <= out_7_7;

         
    when b"101000000" =>reg_data_out <= slv_reg320;     when b"101000001" =>reg_data_out <= slv_reg321;    
    when b"101000010" =>reg_data_out <= slv_reg322;     when b"101000011" =>reg_data_out <= slv_reg323;    
    when b"101000100" =>reg_data_out <= slv_reg324;     when b"101000101" =>reg_data_out <= slv_reg325;    
    when b"101000110" =>reg_data_out <= slv_reg326;     when b"101000111" =>reg_data_out <= slv_reg327;    
    when b"101001000" =>reg_data_out <= slv_reg328;     when b"101001001" =>reg_data_out <= slv_reg329;    
    when b"101001010" =>reg_data_out <= slv_reg330;     when b"101001011" =>reg_data_out <= slv_reg331;    
    when b"101001100" =>reg_data_out <= slv_reg332;     when b"101001101" =>reg_data_out <= slv_reg333;    
    when b"101001110" =>reg_data_out <= slv_reg334;     when b"101001111" =>reg_data_out <= slv_reg335;    
    when b"101010000" =>reg_data_out <= slv_reg336;     when b"101010001" =>reg_data_out <= slv_reg337;    
    when b"101010010" =>reg_data_out <= slv_reg338;     when b"101010011" =>reg_data_out <= slv_reg339;    
    when b"101010100" =>reg_data_out <= slv_reg340;     when b"101010101" =>reg_data_out <= slv_reg341;    
    when b"101010110" =>reg_data_out <= slv_reg342;     when b"101010111" =>reg_data_out <= slv_reg343;    
    when b"101011000" =>reg_data_out <= slv_reg344;     when b"101011001" =>reg_data_out <= slv_reg345;    
    when b"101011010" =>reg_data_out <= slv_reg346;     when b"101011011" =>reg_data_out <= slv_reg347;    
    when b"101011100" =>reg_data_out <= slv_reg348;     when b"101011101" =>reg_data_out <= slv_reg349;    
    when b"101011110" =>reg_data_out <= slv_reg350;     when b"101011111" =>reg_data_out <= slv_reg351;    
    when b"101100000" =>reg_data_out <= slv_reg352;     when b"101100001" =>reg_data_out <= slv_reg353;    
    when b"101100010" =>reg_data_out <= slv_reg354;     when b"101100011" =>reg_data_out <= slv_reg355;    
    when b"101100100" =>reg_data_out <= slv_reg356;     when b"101100101" =>reg_data_out <= slv_reg357;    
    when b"101100110" =>reg_data_out <= slv_reg358;     when b"101100111" =>reg_data_out <= slv_reg359;    
    when b"101101000" =>reg_data_out <= slv_reg360;     when b"101101001" =>reg_data_out <= slv_reg361;    
    when b"101101010" =>reg_data_out <= slv_reg362;     when b"101101011" =>reg_data_out <= slv_reg363;    
    when b"101101100" =>reg_data_out <= slv_reg364;     when b"101101101" =>reg_data_out <= slv_reg365;    
    when b"101101110" =>reg_data_out <= slv_reg366;     when b"101101111" =>reg_data_out <= slv_reg367;    
    when b"101110000" =>reg_data_out <= slv_reg368;     when b"101110001" =>reg_data_out <= slv_reg369;    
    when b"101110010" =>reg_data_out <= slv_reg370;     when b"101110011" =>reg_data_out <= slv_reg371;    
    when b"101110100" =>reg_data_out <= slv_reg372;     when b"101110101" =>reg_data_out <= slv_reg373;    
    when b"101110110" =>reg_data_out <= slv_reg374;     when b"101110111" =>reg_data_out <= slv_reg375;    
    when b"101111000" =>reg_data_out <= slv_reg376;     when b"101111001" =>reg_data_out <= slv_reg377;    
    when b"101111010" =>reg_data_out <= slv_reg378;     when b"101111011" =>reg_data_out <= slv_reg379;    
    when b"101111100" =>reg_data_out <= slv_reg380;     when b"101111101" =>reg_data_out <= slv_reg381;    
    when b"101111110" =>reg_data_out <= slv_reg382;     when b"101111111" =>reg_data_out <= slv_reg383;    
    when b"110000000" =>reg_data_out <= slv_reg384;     when b"110000001" =>reg_data_out <= slv_reg385;    
    when b"110000010" =>reg_data_out <= slv_reg386;     when b"110000011" =>reg_data_out <= slv_reg387;    
    when b"110000100" =>reg_data_out <= slv_reg388;     when b"110000101" =>reg_data_out <= slv_reg389;    
    when b"110000110" =>reg_data_out <= slv_reg390;     when b"110000111" =>reg_data_out <= slv_reg391;    
    when b"110001000" =>reg_data_out <= slv_reg392;     when b"110001001" =>reg_data_out <= slv_reg393;    
    when b"110001010" =>reg_data_out <= slv_reg394;     when b"110001011" =>reg_data_out <= slv_reg395;    
    when b"110001100" =>reg_data_out <= slv_reg396;     when b"110001101" =>reg_data_out <= slv_reg397;    
    when b"110001110" =>reg_data_out <= slv_reg398;     when b"110001111" =>reg_data_out <= slv_reg399;    
    when b"110010000" =>reg_data_out <= slv_reg400;     when b"110010001" =>reg_data_out <= slv_reg401;    
    when b"110010010" =>reg_data_out <= slv_reg402;     when b"110010011" =>reg_data_out <= slv_reg403;    
    when b"110010100" =>reg_data_out <= slv_reg404;     when b"110010101" =>reg_data_out <= slv_reg405;    
    when b"110010110" =>reg_data_out <= slv_reg406;     when b"110010111" =>reg_data_out <= slv_reg407;    
    when b"110011000" =>reg_data_out <= slv_reg408;     when b"110011001" =>reg_data_out <= slv_reg409;    
    when b"110011010" =>reg_data_out <= slv_reg410;     when b"110011011" =>reg_data_out <= slv_reg411;    
    when b"110011100" =>reg_data_out <= slv_reg412;     when b"110011101" =>reg_data_out <= slv_reg413;    
    when b"110011110" =>reg_data_out <= slv_reg414;     when b"110011111" =>reg_data_out <= slv_reg415;    
    when b"110100000" =>reg_data_out <= slv_reg416;     when b"110100001" =>reg_data_out <= slv_reg417;    
    when b"110100010" =>reg_data_out <= slv_reg418;     when b"110100011" =>reg_data_out <= slv_reg419;    
    when b"110100100" =>reg_data_out <= slv_reg420;     when b"110100101" =>reg_data_out <= slv_reg421;    
    when b"110100110" =>reg_data_out <= slv_reg422;     when b"110100111" =>reg_data_out <= slv_reg423;    
    when b"110101000" =>reg_data_out <= slv_reg424;     when b"110101001" =>reg_data_out <= slv_reg425;    
    when b"110101010" =>reg_data_out <= slv_reg426;     when b"110101011" =>reg_data_out <= slv_reg427;    
    when b"110101100" =>reg_data_out <= slv_reg428;     when b"110101101" =>reg_data_out <= slv_reg429;    
    when b"110101110" =>reg_data_out <= slv_reg430;     when b"110101111" =>reg_data_out <= slv_reg431;    
    when b"110110000" =>reg_data_out <= slv_reg432;     when b"110110001" =>reg_data_out <= slv_reg433;    
    when b"110110010" =>reg_data_out <= slv_reg434;     when b"110110011" =>reg_data_out <= slv_reg435;    
    when b"110110100" =>reg_data_out <= slv_reg436;     when b"110110101" =>reg_data_out <= slv_reg437;    
    when b"110110110" =>reg_data_out <= slv_reg438;     when b"110110111" =>reg_data_out <= slv_reg439;    
    when b"110111000" =>reg_data_out <= slv_reg440;     when b"110111001" =>reg_data_out <= slv_reg441;    
    when b"110111010" =>reg_data_out <= slv_reg442;     when b"110111011" =>reg_data_out <= slv_reg443;    
    when b"110111100" =>reg_data_out <= slv_reg444;     when b"110111101" =>reg_data_out <= slv_reg445;    
    when b"110111110" =>reg_data_out <= slv_reg446;     when b"110111111" =>reg_data_out <= slv_reg447;    
    when b"111000000" =>reg_data_out <= slv_reg448;     when b"111000001" =>reg_data_out <= slv_reg449;    
    when b"111000010" =>reg_data_out <= slv_reg450;     when b"111000011" =>reg_data_out <= slv_reg451; 
    when b"111000100" =>reg_data_out <= slv_reg452;     when b"111000101" =>reg_data_out <= slv_reg453;    
    when b"111000110" =>reg_data_out <= slv_reg454;     when b"111000111" =>reg_data_out <= slv_reg455;    
    when b"111001000" =>reg_data_out <= slv_reg456;     when b"111001001" =>reg_data_out <= slv_reg457;    
    when b"111001010" =>reg_data_out <= slv_reg458;     when b"111001011" =>reg_data_out <= slv_reg459;    
    when b"111001100" =>reg_data_out <= slv_reg460;     when b"111001101" =>reg_data_out <= slv_reg461;    
    when b"111001110" =>reg_data_out <= slv_reg462;     when b"111001111" =>reg_data_out <= slv_reg463;    
    when b"111010000" =>reg_data_out <= slv_reg464;     when b"111010001" =>reg_data_out <= slv_reg465;    
    when b"111010010" =>reg_data_out <= slv_reg466;     when b"111010011" =>reg_data_out <= slv_reg467;    
    when b"111010100" =>reg_data_out <= slv_reg468;     when b"111010101" =>reg_data_out <= slv_reg469;    
    when b"111010110" =>reg_data_out <= slv_reg470;     when b"111010111" =>reg_data_out <= slv_reg471;    
    when b"111011000" =>reg_data_out <= slv_reg472;     when b"111011001" =>reg_data_out <= slv_reg473;    
    when b"111011010" =>reg_data_out <= slv_reg474;     when b"111011011" =>reg_data_out <= slv_reg475;    
    when b"111011100" =>reg_data_out <= slv_reg476;     when b"111011101" =>reg_data_out <= slv_reg477;    
    when b"111011110" =>reg_data_out <= slv_reg478;     when b"111011111" =>reg_data_out <= slv_reg479;    
    when b"111100000" =>reg_data_out <= slv_reg480;     when b"111100001" =>reg_data_out <= slv_reg481;    
    when b"111100010" =>reg_data_out <= slv_reg482;     when b"111100011" =>reg_data_out <= slv_reg483;    
    when b"111100100" =>reg_data_out <= slv_reg484;     when b"111100101" =>reg_data_out <= slv_reg485;    
    when b"111100110" =>reg_data_out <= slv_reg486;     when b"111100111" =>reg_data_out <= slv_reg487;    
    when b"111101000" =>reg_data_out <= slv_reg488;     when b"111101001" =>reg_data_out <= slv_reg489;    
    when b"111101010" =>reg_data_out <= slv_reg490;     when b"111101011" =>reg_data_out <= slv_reg491;    
    when b"111101100" =>reg_data_out <= slv_reg492;     when b"111101101" =>reg_data_out <= slv_reg493;    
    when b"111101110" =>reg_data_out <= slv_reg494;     when b"111101111" =>reg_data_out <= slv_reg495;    
    when b"111110000" =>reg_data_out <= slv_reg496;     when b"111110001" =>reg_data_out <= slv_reg497;    
    when b"111110010" =>reg_data_out <= slv_reg498;     when b"111110011" =>reg_data_out <= slv_reg499;    
    when b"111110100" =>reg_data_out <= slv_reg500;     when b"111110101" =>reg_data_out <= slv_reg501;    
    when b"111110110" =>reg_data_out <= slv_reg502;     when b"111110111" =>reg_data_out <= slv_reg503;    
    when b"111111000" =>reg_data_out <= slv_reg504;     when b"111111001" =>reg_data_out <= slv_reg505;    
    when b"111111010" =>reg_data_out <= slv_reg506;     when b"111111011" =>reg_data_out <= slv_reg507;    
    when b"111111100" =>reg_data_out <= slv_reg508;     when b"111111101" =>reg_data_out <= slv_reg509;    
    when b"111111110" =>reg_data_out <= slv_reg510;     when b"111111111" =>reg_data_out <= slv_reg511;
--  = # = # = # = # = # = # = # = # = # = # = # = # = # = # = # = # = # = # = # = # = # = # = # = # = # = # = # = #
    
    when others =>reg_data_out  <= (others => '0');
    end case;
end process; 



	
--  = # = # = # = # = # = # = # = # = # = # = # = # = # = # = # = # = # = # = # = # = # = # = # = # = # = # = # = # 
--  = # = # = # = # = # = # = # = # = # = # = # = # = # = # = # = # = # = # = # = # = # = # = # = # = # = # = # = #

    
--  = # = # = # = # = # = # = # = # = # = # = # = # = # = # = # = # = # = # = # = # = # = # = # = # = # = # = # = #
--  = # = # = # = # = # = # = # = # = # = # = # = # = # = # = # = # = # = # = # = # = # = # = # = # = # = # = # = #


--  S T O P             S T O P             S T O P             S T O P             S T O P             S T O P

--          H E R E             H E R E             H E R E             H E R E             H E R E             H E R E


	
--  = # = # = # = # = # = # = # = # = # = # = # = # = # = # = # = # = # = # = # = # = # = # = # = # = # = # = # = # 
--  = # = # = # = # = # = # = # = # = # = # = # = # = # = # = # = # = # = # = # = # = # = # = # = # = # = # = # = #

    
--  = # = # = # = # = # = # = # = # = # = # = # = # = # = # = # = # = # = # = # = # = # = # = # = # = # = # = # = #
--  = # = # = # = # = # = # = # = # = # = # = # = # = # = # = # = # = # = # = # = # = # = # = # = # = # = # = # = #



	S_AXI_AWREADY  <= axi_awready;
	S_AXI_WREADY   <= axi_wready;
	S_AXI_BRESP	   <= axi_bresp;
	S_AXI_BVALID   <= axi_bvalid;
	S_AXI_ARREADY  <= axi_arready;
	S_AXI_RDATA    <= axi_rdata;
	S_AXI_RRESP    <= axi_rresp;
	S_AXI_RVALID   <= axi_rvalid;
	

	process (S_AXI_ACLK)
	begin
	  if rising_edge(S_AXI_ACLK) then 
	    if S_AXI_ARESETN = '0' then
	      axi_awready <= '0';
	      aw_en <= '1';
	    else
	      if (axi_awready = '0' and S_AXI_AWVALID = '1' and S_AXI_WVALID = '1' and aw_en = '1') then
	        axi_awready <= '1';
	        elsif (S_AXI_BREADY = '1' and axi_bvalid = '1') then
	            aw_en <= '1';
	        	axi_awready <= '0';
	      else
	        axi_awready <= '0';
	      end if;
	    end if;
	  end if;
	end process;

	process (S_AXI_ACLK)
	begin
	  if rising_edge(S_AXI_ACLK) then 
	    if S_AXI_ARESETN = '0' then
	      axi_awaddr <= (others => '0');
	    else
	      if (axi_awready = '0' and S_AXI_AWVALID = '1' and S_AXI_WVALID = '1' and aw_en = '1') then
	        axi_awaddr <= S_AXI_AWADDR;
	      end if;
	    end if;
	  end if;                   
	end process; 

	process (S_AXI_ACLK)
	begin
	  if rising_edge(S_AXI_ACLK) then 
	    if S_AXI_ARESETN = '0' then
	      axi_wready <= '0';
	    else
	      if (axi_wready = '0' and S_AXI_WVALID = '1' and S_AXI_AWVALID = '1' and aw_en = '1') then
	        axi_wready <= '1';
	      else
	        axi_wready <= '0';
	      end if;
	    end if;
	  end if;
	end process; 

	--RESET
	slv_reg_wren <= axi_wready and S_AXI_WVALID and axi_awready and S_AXI_AWVALID ;
    
    


	process (S_AXI_ACLK)
	variable loc_addr :std_logic_vector(OPT_MEM_ADDR_BITS downto 0); 
	begin
	  if rising_edge(S_AXI_ACLK) then 
	    if S_AXI_ARESETN = '0' then
            slv_reg0<=(others=>'0');   slv_reg1<=(others=>'0');   slv_reg2<=(others=>'0');   slv_reg3<=(others=>'0'); 
            slv_reg4<=(others=>'0');   slv_reg5<=(others=>'0');   slv_reg6<=(others=>'0');   slv_reg7<=(others=>'0'); 
            slv_reg8<=(others=>'0');   slv_reg9<=(others=>'0');   slv_reg10<=(others=>'0');  slv_reg11<=(others=>'0'); 
            slv_reg12<=(others=>'0');  slv_reg13<=(others=>'0');  slv_reg14<=(others=>'0');  slv_reg15<=(others=>'0'); 
            slv_reg16<=(others=>'0');  slv_reg17<=(others=>'0');  slv_reg18<=(others=>'0');  slv_reg19<=(others=>'0'); 
            slv_reg20<=(others=>'0');  slv_reg21<=(others=>'0');  slv_reg22<=(others=>'0');  slv_reg23<=(others=>'0'); 
            slv_reg24<=(others=>'0');  slv_reg25<=(others=>'0');  slv_reg26<=(others=>'0');  slv_reg27<=(others=>'0'); 
            slv_reg28<=(others=>'0');  slv_reg29<=(others=>'0');  slv_reg30<=(others=>'0');  slv_reg31<=(others=>'0'); 
            slv_reg32<=(others=>'0');  slv_reg33<=(others=>'0');  slv_reg34<=(others=>'0');  slv_reg35<=(others=>'0'); 
            slv_reg36<=(others=>'0');  slv_reg37<=(others=>'0');  slv_reg38<=(others=>'0');  slv_reg39<=(others=>'0'); 
            slv_reg40<=(others=>'0');  slv_reg41<=(others=>'0');  slv_reg42<=(others=>'0');  slv_reg43<=(others=>'0'); 
            slv_reg44<=(others=>'0');  slv_reg45<=(others=>'0');  slv_reg46<=(others=>'0');  slv_reg47<=(others=>'0'); 
            slv_reg48<=(others=>'0');  slv_reg49<=(others=>'0');  slv_reg50<=(others=>'0');  slv_reg51<=(others=>'0'); 
            slv_reg52<=(others=>'0');  slv_reg53<=(others=>'0');  slv_reg54<=(others=>'0');  slv_reg55<=(others=>'0'); 
            slv_reg56<=(others=>'0');  slv_reg57<=(others=>'0');  slv_reg58<=(others=>'0');  slv_reg59<=(others=>'0'); 
            slv_reg60<=(others=>'0');  slv_reg61<=(others=>'0');  slv_reg62<=(others=>'0');  slv_reg63<=(others=>'0');
             
            slv_reg64<=(others=>'0');  slv_reg65<=(others=>'0');  slv_reg66<=(others=>'0');  slv_reg67<=(others=>'0'); 
            slv_reg68<=(others=>'0');  slv_reg69<=(others=>'0');  slv_reg70<=(others=>'0');  slv_reg71<=(others=>'0'); 
            slv_reg72<=(others=>'0');  slv_reg73<=(others=>'0');  slv_reg74<=(others=>'0');  slv_reg75<=(others=>'0'); 
            slv_reg76<=(others=>'0');  slv_reg77<=(others=>'0');  slv_reg78<=(others=>'0');  slv_reg79<=(others=>'0'); 
            slv_reg80<=(others=>'0');  slv_reg81<=(others=>'0');  slv_reg82<=(others=>'0');  slv_reg83<=(others=>'0'); 
            slv_reg84<=(others=>'0');  slv_reg85<=(others=>'0');  slv_reg86<=(others=>'0');  slv_reg87<=(others=>'0'); 
            slv_reg88<=(others=>'0');  slv_reg89<=(others=>'0');  slv_reg90<=(others=>'0');  slv_reg91<=(others=>'0'); 
            slv_reg92<=(others=>'0');  slv_reg93<=(others=>'0');  slv_reg94<=(others=>'0');  slv_reg95<=(others=>'0'); 
            slv_reg96<=(others=>'0');  slv_reg97<=(others=>'0');  slv_reg98<=(others=>'0');  slv_reg99<=(others=>'0');
            slv_reg100<=(others=>'0'); slv_reg101<=(others=>'0'); slv_reg102<=(others=>'0'); slv_reg103<=(others=>'0'); 
            slv_reg104<=(others=>'0'); slv_reg105<=(others=>'0'); slv_reg106<=(others=>'0'); slv_reg107<=(others=>'0'); 
            slv_reg108<=(others=>'0'); slv_reg109<=(others=>'0'); slv_reg110<=(others=>'0'); slv_reg111<=(others=>'0'); 
            slv_reg112<=(others=>'0'); slv_reg113<=(others=>'0'); slv_reg114<=(others=>'0'); slv_reg115<=(others=>'0'); 
            slv_reg116<=(others=>'0'); slv_reg117<=(others=>'0'); slv_reg118<=(others=>'0'); slv_reg119<=(others=>'0'); 
            slv_reg120<=(others=>'0'); slv_reg121<=(others=>'0'); slv_reg122<=(others=>'0'); slv_reg123<=(others=>'0'); 
            slv_reg124<=(others=>'0'); slv_reg125<=(others=>'0'); slv_reg126<=(others=>'0'); slv_reg127<=(others=>'0');
             
            slv_reg128<=(others=>'0'); slv_reg129<=(others=>'0'); slv_reg130<=(others=>'0'); slv_reg131<=(others=>'0'); 
            slv_reg132<=(others=>'0'); slv_reg133<=(others=>'0'); slv_reg134<=(others=>'0'); slv_reg135<=(others=>'0'); 
            slv_reg136<=(others=>'0'); slv_reg137<=(others=>'0'); slv_reg138<=(others=>'0'); slv_reg139<=(others=>'0');
            slv_reg140<=(others=>'0'); slv_reg141<=(others=>'0'); slv_reg142<=(others=>'0'); slv_reg143<=(others=>'0'); 
            slv_reg144<=(others=>'0'); slv_reg145<=(others=>'0'); slv_reg146<=(others=>'0'); slv_reg147<=(others=>'0'); 
            slv_reg148<=(others=>'0'); slv_reg149<=(others=>'0'); slv_reg150<=(others=>'0'); slv_reg151<=(others=>'0'); 
            slv_reg152<=(others=>'0'); slv_reg153<=(others=>'0'); slv_reg154<=(others=>'0'); slv_reg155<=(others=>'0'); 
            slv_reg156<=(others=>'0'); slv_reg157<=(others=>'0'); slv_reg158<=(others=>'0'); slv_reg159<=(others=>'0');
            slv_reg160<=(others=>'0'); slv_reg161<=(others=>'0'); slv_reg162<=(others=>'0'); slv_reg163<=(others=>'0'); 
            slv_reg164<=(others=>'0'); slv_reg165<=(others=>'0'); slv_reg166<=(others=>'0'); slv_reg167<=(others=>'0'); 
            slv_reg168<=(others=>'0'); slv_reg169<=(others=>'0'); slv_reg170<=(others=>'0'); slv_reg171<=(others=>'0'); 
            slv_reg172<=(others=>'0'); slv_reg173<=(others=>'0'); slv_reg174<=(others=>'0'); slv_reg175<=(others=>'0'); 
            slv_reg176<=(others=>'0'); slv_reg177<=(others=>'0'); slv_reg178<=(others=>'0'); slv_reg179<=(others=>'0'); 
            slv_reg180<=(others=>'0'); slv_reg181<=(others=>'0'); slv_reg182<=(others=>'0'); slv_reg183<=(others=>'0'); 
            slv_reg184<=(others=>'0'); slv_reg185<=(others=>'0'); slv_reg186<=(others=>'0'); slv_reg187<=(others=>'0'); 
            slv_reg188<=(others=>'0'); slv_reg189<=(others=>'0'); slv_reg190<=(others=>'0'); slv_reg191<=(others=>'0'); 
            
            slv_reg192<=(others=>'0'); slv_reg193<=(others=>'0'); slv_reg194<=(others=>'0'); slv_reg195<=(others=>'0'); 
            slv_reg196<=(others=>'0'); slv_reg197<=(others=>'0'); slv_reg198<=(others=>'0'); slv_reg199<=(others=>'0'); 
            slv_reg200<=(others=>'0'); slv_reg201<=(others=>'0'); slv_reg202<=(others=>'0'); slv_reg203<=(others=>'0'); 
            slv_reg204<=(others=>'0'); slv_reg205<=(others=>'0'); slv_reg206<=(others=>'0'); slv_reg207<=(others=>'0'); 
            slv_reg208<=(others=>'0'); slv_reg209<=(others=>'0'); slv_reg210<=(others=>'0'); slv_reg211<=(others=>'0'); 
            slv_reg212<=(others=>'0'); slv_reg213<=(others=>'0'); slv_reg214<=(others=>'0'); slv_reg215<=(others=>'0'); 
            slv_reg216<=(others=>'0'); slv_reg217<=(others=>'0'); slv_reg218<=(others=>'0'); slv_reg219<=(others=>'0'); 
            slv_reg220<=(others=>'0'); slv_reg221<=(others=>'0'); slv_reg222<=(others=>'0'); slv_reg223<=(others=>'0'); 
            slv_reg224<=(others=>'0'); slv_reg225<=(others=>'0'); slv_reg226<=(others=>'0'); slv_reg227<=(others=>'0'); 
            slv_reg228<=(others=>'0'); slv_reg229<=(others=>'0'); slv_reg230<=(others=>'0'); slv_reg231<=(others=>'0'); 
            slv_reg232<=(others=>'0'); slv_reg233<=(others=>'0'); slv_reg234<=(others=>'0'); slv_reg235<=(others=>'0'); 
            slv_reg236<=(others=>'0'); slv_reg237<=(others=>'0'); slv_reg238<=(others=>'0'); slv_reg239<=(others=>'0'); 
            slv_reg240<=(others=>'0'); slv_reg241<=(others=>'0'); slv_reg242<=(others=>'0'); slv_reg243<=(others=>'0'); 
            slv_reg244<=(others=>'0'); slv_reg245<=(others=>'0'); slv_reg246<=(others=>'0'); slv_reg247<=(others=>'0'); 
            slv_reg248<=(others=>'0'); slv_reg249<=(others=>'0'); slv_reg250<=(others=>'0'); slv_reg251<=(others=>'0'); 
            slv_reg252<=(others=>'0'); slv_reg253<=(others=>'0'); slv_reg254<=(others=>'0'); slv_reg255<=(others=>'0');
             
            slv_reg256<=(others=>'0'); slv_reg257<=(others=>'0'); slv_reg258<=(others=>'0'); slv_reg259<=(others=>'0'); 
            slv_reg260<=(others=>'0'); slv_reg261<=(others=>'0'); slv_reg262<=(others=>'0'); slv_reg263<=(others=>'0'); 
            slv_reg264<=(others=>'0'); slv_reg265<=(others=>'0'); slv_reg266<=(others=>'0'); slv_reg267<=(others=>'0'); 
            slv_reg268<=(others=>'0'); slv_reg269<=(others=>'0'); slv_reg270<=(others=>'0'); slv_reg271<=(others=>'0'); 
            slv_reg272<=(others=>'0'); slv_reg273<=(others=>'0'); slv_reg274<=(others=>'0'); slv_reg275<=(others=>'0'); 
            slv_reg276<=(others=>'0'); slv_reg277<=(others=>'0'); slv_reg278<=(others=>'0'); slv_reg279<=(others=>'0'); 
            slv_reg280<=(others=>'0'); slv_reg281<=(others=>'0'); slv_reg282<=(others=>'0'); slv_reg283<=(others=>'0'); 
            slv_reg284<=(others=>'0'); slv_reg285<=(others=>'0'); slv_reg286<=(others=>'0'); slv_reg287<=(others=>'0'); 
            slv_reg288<=(others=>'0'); slv_reg289<=(others=>'0'); slv_reg290<=(others=>'0'); slv_reg291<=(others=>'0'); 
            slv_reg292<=(others=>'0'); slv_reg293<=(others=>'0'); slv_reg294<=(others=>'0'); slv_reg295<=(others=>'0'); 
            slv_reg296<=(others=>'0'); slv_reg297<=(others=>'0'); slv_reg298<=(others=>'0'); slv_reg299<=(others=>'0'); 
            slv_reg300<=(others=>'0'); slv_reg301<=(others=>'0'); slv_reg302<=(others=>'0'); slv_reg303<=(others=>'0'); 
            slv_reg304<=(others=>'0'); slv_reg305<=(others=>'0'); slv_reg306<=(others=>'0'); slv_reg307<=(others=>'0'); 
            slv_reg308<=(others=>'0'); slv_reg309<=(others=>'0'); slv_reg310<=(others=>'0'); slv_reg311<=(others=>'0'); 
            slv_reg312<=(others=>'0'); slv_reg313<=(others=>'0'); slv_reg314<=(others=>'0'); slv_reg315<=(others=>'0'); 
            slv_reg316<=(others=>'0'); slv_reg317<=(others=>'0'); slv_reg318<=(others=>'0'); slv_reg319<=(others=>'0');
             
            slv_reg320<=(others=>'0'); slv_reg321<=(others=>'0'); slv_reg322<=(others=>'0'); slv_reg323<=(others=>'0'); 
            slv_reg324<=(others=>'0'); slv_reg325<=(others=>'0'); slv_reg326<=(others=>'0'); slv_reg327<=(others=>'0'); 
            slv_reg328<=(others=>'0'); slv_reg329<=(others=>'0'); slv_reg330<=(others=>'0'); slv_reg331<=(others=>'0'); 
            slv_reg332<=(others=>'0'); slv_reg333<=(others=>'0'); slv_reg334<=(others=>'0'); slv_reg335<=(others=>'0'); 
            slv_reg336<=(others=>'0'); slv_reg337<=(others=>'0'); slv_reg338<=(others=>'0'); slv_reg339<=(others=>'0'); 
            slv_reg340<=(others=>'0'); slv_reg341<=(others=>'0'); slv_reg342<=(others=>'0'); slv_reg343<=(others=>'0'); 
            slv_reg344<=(others=>'0'); slv_reg345<=(others=>'0'); slv_reg346<=(others=>'0'); slv_reg347<=(others=>'0'); 
            slv_reg348<=(others=>'0'); slv_reg349<=(others=>'0'); slv_reg350<=(others=>'0'); slv_reg351<=(others=>'0'); 
            slv_reg352<=(others=>'0'); slv_reg353<=(others=>'0'); slv_reg354<=(others=>'0'); slv_reg355<=(others=>'0'); 
            slv_reg356<=(others=>'0'); slv_reg357<=(others=>'0'); slv_reg358<=(others=>'0'); slv_reg359<=(others=>'0'); 
            slv_reg360<=(others=>'0'); slv_reg361<=(others=>'0'); slv_reg362<=(others=>'0'); slv_reg363<=(others=>'0'); 
            slv_reg364<=(others=>'0'); slv_reg365<=(others=>'0'); slv_reg366<=(others=>'0'); slv_reg367<=(others=>'0'); 
            slv_reg368<=(others=>'0'); slv_reg369<=(others=>'0'); slv_reg370<=(others=>'0'); slv_reg371<=(others=>'0'); 
            slv_reg372<=(others=>'0'); slv_reg373<=(others=>'0'); slv_reg374<=(others=>'0'); slv_reg375<=(others=>'0'); 
            slv_reg376<=(others=>'0'); slv_reg377<=(others=>'0'); slv_reg378<=(others=>'0'); slv_reg379<=(others=>'0'); 
            slv_reg380<=(others=>'0'); slv_reg381<=(others=>'0'); slv_reg382<=(others=>'0'); slv_reg383<=(others=>'0');
             
            slv_reg384<=(others=>'0'); slv_reg385<=(others=>'0'); slv_reg386<=(others=>'0'); slv_reg387<=(others=>'0'); 
            slv_reg388<=(others=>'0'); slv_reg389<=(others=>'0'); slv_reg390<=(others=>'0'); slv_reg391<=(others=>'0'); 
            slv_reg392<=(others=>'0'); slv_reg393<=(others=>'0'); slv_reg394<=(others=>'0'); slv_reg395<=(others=>'0'); 
            slv_reg396<=(others=>'0'); slv_reg397<=(others=>'0'); slv_reg398<=(others=>'0'); slv_reg399<=(others=>'0'); 
            slv_reg400<=(others=>'0'); slv_reg401<=(others=>'0'); slv_reg402<=(others=>'0'); slv_reg403<=(others=>'0'); 
            slv_reg404<=(others=>'0'); slv_reg405<=(others=>'0'); slv_reg406<=(others=>'0'); slv_reg407<=(others=>'0'); 
            slv_reg408<=(others=>'0'); slv_reg409<=(others=>'0'); slv_reg410<=(others=>'0'); slv_reg411<=(others=>'0'); 
            slv_reg412<=(others=>'0'); slv_reg413<=(others=>'0'); slv_reg414<=(others=>'0'); slv_reg415<=(others=>'0'); 
            slv_reg416<=(others=>'0'); slv_reg417<=(others=>'0'); slv_reg418<=(others=>'0'); slv_reg419<=(others=>'0'); 
            slv_reg420<=(others=>'0'); slv_reg421<=(others=>'0'); slv_reg422<=(others=>'0'); slv_reg423<=(others=>'0'); 
            slv_reg424<=(others=>'0'); slv_reg425<=(others=>'0'); slv_reg426<=(others=>'0'); slv_reg427<=(others=>'0'); 
            slv_reg428<=(others=>'0'); slv_reg429<=(others=>'0'); slv_reg430<=(others=>'0'); slv_reg431<=(others=>'0'); 
            slv_reg432<=(others=>'0'); slv_reg433<=(others=>'0'); slv_reg434<=(others=>'0'); slv_reg435<=(others=>'0'); 
            slv_reg436<=(others=>'0'); slv_reg437<=(others=>'0'); slv_reg438<=(others=>'0'); slv_reg439<=(others=>'0'); 
            slv_reg440<=(others=>'0'); slv_reg441<=(others=>'0'); slv_reg442<=(others=>'0'); slv_reg443<=(others=>'0'); 
            slv_reg444<=(others=>'0'); slv_reg445<=(others=>'0'); slv_reg446<=(others=>'0'); slv_reg447<=(others=>'0');
             
            slv_reg448<=(others=>'0'); slv_reg449<=(others=>'0'); slv_reg450<=(others=>'0'); slv_reg451<=(others=>'0'); 
            slv_reg452<=(others=>'0'); slv_reg453<=(others=>'0'); slv_reg454<=(others=>'0'); slv_reg455<=(others=>'0'); 
            slv_reg456<=(others=>'0'); slv_reg457<=(others=>'0'); slv_reg458<=(others=>'0'); slv_reg459<=(others=>'0'); 
            slv_reg460<=(others=>'0'); slv_reg461<=(others=>'0'); slv_reg462<=(others=>'0'); slv_reg463<=(others=>'0'); 
            slv_reg464<=(others=>'0'); slv_reg465<=(others=>'0'); slv_reg466<=(others=>'0'); slv_reg467<=(others=>'0'); 
            slv_reg468<=(others=>'0'); slv_reg469<=(others=>'0'); slv_reg470<=(others=>'0'); slv_reg471<=(others=>'0'); 
            slv_reg472<=(others=>'0'); slv_reg473<=(others=>'0'); slv_reg474<=(others=>'0'); slv_reg475<=(others=>'0'); 
            slv_reg476<=(others=>'0'); slv_reg477<=(others=>'0'); slv_reg478<=(others=>'0'); slv_reg479<=(others=>'0'); 
            slv_reg480<=(others=>'0'); slv_reg481<=(others=>'0'); slv_reg482<=(others=>'0'); slv_reg483<=(others=>'0'); 
            slv_reg484<=(others=>'0'); slv_reg485<=(others=>'0'); slv_reg486<=(others=>'0'); slv_reg487<=(others=>'0'); 
            slv_reg488<=(others=>'0'); slv_reg489<=(others=>'0'); slv_reg490<=(others=>'0'); slv_reg491<=(others=>'0'); 
            slv_reg492<=(others=>'0'); slv_reg493<=(others=>'0'); slv_reg494<=(others=>'0'); slv_reg495<=(others=>'0'); 
            slv_reg496<=(others=>'0'); slv_reg497<=(others=>'0'); slv_reg498<=(others=>'0'); slv_reg499<=(others=>'0'); 
            slv_reg500<=(others=>'0'); slv_reg501<=(others=>'0'); slv_reg502<=(others=>'0'); slv_reg503<=(others=>'0'); 
            slv_reg504<=(others=>'0'); slv_reg505<=(others=>'0'); slv_reg506<=(others=>'0'); slv_reg507<=(others=>'0'); 
            slv_reg508<=(others=>'0'); slv_reg509<=(others=>'0'); slv_reg510<=(others=>'0'); slv_reg511<=(others=>'0');     
	else
	  loc_addr := axi_awaddr(ADDR_LSB + OPT_MEM_ADDR_BITS downto ADDR_LSB);
	  if (slv_reg_wren = '1') then
	
        case loc_addr is
           when b"000000000" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg0(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;        end loop;
           when b"000000001" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg1(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;        end loop;
           when b"000000010" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg2(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;        end loop;
           when b"000000011" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg3(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;        end loop;
           when b"000000100" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg4(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;        end loop;
           when b"000000101" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg5(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;        end loop;
           when b"000000110" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg6(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;        end loop;
           when b"000000111" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg7(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;        end loop;
           when b"000001000" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg8(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;        end loop;
           when b"000001001" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg9(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;        end loop;
           when b"000001010" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg10(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;        end loop;
           when b"000001011" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg11(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;        end loop;
           when b"000001100" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg12(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;        end loop;
           when b"000001101" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg13(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;        end loop;
           when b"000001110" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg14(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;        end loop;
           when b"000001111" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg15(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;        end loop;
           when b"000010000" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg16(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;        end loop;
           when b"000010001" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg17(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;        end loop;
           when b"000010010" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg18(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;        end loop;
           when b"000010011" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg19(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;        end loop;
           when b"000010100" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg20(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;        end loop;
           when b"000010101" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg21(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;        end loop;
           when b"000010110" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg22(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;        end loop;
           when b"000010111" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg23(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;        end loop;
           when b"000011000" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg24(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;        end loop;
           when b"000011001" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg25(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;        end loop;
           when b"000011010" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg26(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;        end loop;
           when b"000011011" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg27(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;        end loop;
           when b"000011100" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg28(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"000011101" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg29(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"000011110" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg30(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"000011111" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg31(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"000100000" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg32(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"000100001" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg33(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"000100010" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg34(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"000100011" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg35(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"000100100" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg36(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"000100101" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg37(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"000100110" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg38(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"000100111" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg39(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"000101000" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg40(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"000101001" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg41(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"000101010" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg42(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"000101011" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg43(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"000101100" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg44(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"000101101" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg45(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"000101110" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg46(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"000101111" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg47(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"000110000" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg48(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"000110001" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg49(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"000110010" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg50(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"000110011" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg51(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"000110100" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg52(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"000110101" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg53(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"000110110" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg54(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"000110111" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg55(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"000111000" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg56(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"000111001" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg57(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"000111010" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg58(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"000111011" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg59(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"000111100" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg60(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"000111101" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg61(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"000111110" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg62(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"000111111" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg63(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"001000000" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg64(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"001000001" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg65(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"001000010" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg66(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"001000011" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg67(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"001000100" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg68(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"001000101" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg69(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"001000110" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg70(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"001000111" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg71(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"001001000" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg72(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"001001001" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg73(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"001001010" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg74(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"001001011" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg75(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"001001100" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg76(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"001001101" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg77(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"001001110" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg78(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"001001111" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg79(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"001010000" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg80(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"001010001" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg81(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"001010010" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg82(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"001010011" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg83(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"001010100" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg84(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"001010101" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg85(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"001010110" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg86(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"001010111" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg87(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"001011000" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg88(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"001011001" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg89(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"001011010" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg90(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"001011011" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg91(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"001011100" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg92(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"001011101" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg93(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"001011110" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg94(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"001011111" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg95(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"001100000" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg96(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"001100001" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg97(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"001100010" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg98(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"001100011" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg99(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"001100100" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg100(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"001100101" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg101(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"001100110" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg102(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"001100111" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg103(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"001101000" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg104(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"001101001" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg105(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"001101010" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg106(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"001101011" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg107(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"001101100" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg108(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"001101101" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg109(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"001101110" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg110(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"001101111" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg111(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"001110000" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg112(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"001110001" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg113(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"001110010" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg114(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"001110011" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg115(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"001110100" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg116(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"001110101" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg117(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"001110110" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg118(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"001110111" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg119(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"001111000" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg120(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"001111001" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg121(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"001111010" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg122(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"001111011" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg123(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"001111100" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg124(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"001111101" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg125(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"001111110" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg126(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"001111111" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg127(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"010000000" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg128(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"010000001" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg129(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"010000010" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg130(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"010000011" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg131(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"010000100" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg132(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"010000101" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg133(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"010000110" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg134(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"010000111" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg135(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"010001000" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg136(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"010001001" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg137(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"010001010" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg138(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"010001011" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg139(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"010001100" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg140(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"010001101" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg141(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"010001110" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg142(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"010001111" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg143(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"010010000" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg144(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"010010001" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg145(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"010010010" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg146(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"010010011" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg147(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"010010100" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg148(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"010010101" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg149(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"010010110" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg150(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"010010111" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg151(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"010011000" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg152(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"010011001" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg153(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"010011010" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg154(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"010011011" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg155(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"010011100" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg156(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"010011101" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg157(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"010011110" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg158(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"010011111" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg159(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"010100000" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg160(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"010100001" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg161(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"010100010" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg162(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"010100011" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg163(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"010100100" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg164(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"010100101" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg165(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"010100110" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg166(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"010100111" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg167(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"010101000" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg168(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"010101001" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg169(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"010101010" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg170(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"010101011" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg171(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"010101100" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg172(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"010101101" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg173(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"010101110" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg174(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"010101111" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg175(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"010110000" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg176(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"010110001" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg177(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"010110010" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg178(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"010110011" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg179(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"010110100" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg180(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"010110101" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg181(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"010110110" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg182(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"010110111" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg183(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"010111000" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg184(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"010111001" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg185(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"010111010" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg186(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"010111011" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg187(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"010111100" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg188(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"010111101" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg189(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"010111110" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg190(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"010111111" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg191(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"011000000" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg192(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"011000001" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg193(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"011000010" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg194(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"011000011" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg195(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"011000100" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg196(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"011000101" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg197(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"011000110" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg198(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"011000111" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg199(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"011001000" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg200(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"011001001" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg201(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"011001010" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg202(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"011001011" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg203(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"011001100" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg204(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"011001101" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg205(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"011001110" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg206(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"011001111" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg207(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"011010000" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg208(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"011010001" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg209(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"011010010" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg210(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"011010011" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg211(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"011010100" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg212(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"011010101" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg213(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"011010110" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg214(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"011010111" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg215(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"011011000" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg216(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"011011001" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg217(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"011011010" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg218(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"011011011" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg219(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"011011100" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg220(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"011011101" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg221(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"011011110" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg222(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"011011111" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg223(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"011100000" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg224(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"011100001" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg225(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"011100010" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg226(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"011100011" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg227(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"011100100" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg228(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"011100101" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg229(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"011100110" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg230(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"011100111" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg231(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"011101000" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg232(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"011101001" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg233(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"011101010" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg234(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"011101011" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg235(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"011101100" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg236(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"011101101" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg237(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"011101110" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg238(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"011101111" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg239(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"011110000" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg240(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"011110001" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg241(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"011110010" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg242(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"011110011" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg243(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"011110100" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg244(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"011110101" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg245(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"011110110" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg246(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"011110111" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg247(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"011111000" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg248(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"011111001" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg249(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"011111010" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg250(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"011111011" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg251(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"011111100" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg252(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"011111101" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg253(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"011111110" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg254(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"011111111" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg255(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"100000000" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg256(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"100000001" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg257(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"100000010" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg258(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"100000011" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg259(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"100000100" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg260(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"100000101" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg261(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"100000110" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg262(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"100000111" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg263(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"100001000" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg264(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"100001001" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg265(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"100001010" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg266(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"100001011" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg267(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"100001100" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg268(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"100001101" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg269(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"100001110" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg270(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"100001111" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg271(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"100010000" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg272(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"100010001" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg273(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"100010010" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg274(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"100010011" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg275(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"100010100" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg276(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"100010101" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg277(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"100010110" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg278(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"100010111" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg279(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"100011000" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg280(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"100011001" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg281(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"100011010" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg282(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"100011011" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg283(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"100011100" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg284(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"100011101" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg285(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"100011110" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg286(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"100011111" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg287(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"100100000" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg288(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"100100001" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg289(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"100100010" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg290(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"100100011" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg291(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"100100100" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg292(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"100100101" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg293(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"100100110" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg294(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"100100111" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg295(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"100101000" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg296(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"100101001" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg297(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"100101010" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg298(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"100101011" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg299(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"100101100" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg300(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"100101101" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg301(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"100101110" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg302(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"100101111" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg303(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"100110000" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg304(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"100110001" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg305(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"100110010" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg306(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"100110011" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg307(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"100110100" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg308(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"100110101" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg309(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"100110110" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg310(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"100110111" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg311(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"100111000" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg312(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"100111001" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg313(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"100111010" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg314(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"100111011" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg315(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"100111100" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg316(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"100111101" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg317(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"100111110" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg318(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"100111111" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg319(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"101000000" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg320(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"101000001" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg321(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"101000010" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg322(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"101000011" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg323(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"101000100" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg324(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"101000101" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg325(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"101000110" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg326(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"101000111" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg327(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"101001000" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg328(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"101001001" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg329(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"101001010" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg330(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"101001011" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg331(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"101001100" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg332(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"101001101" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg333(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"101001110" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg334(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"101001111" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg335(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"101010000" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg336(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"101010001" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg337(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"101010010" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg338(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"101010011" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg339(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"101010100" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg340(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"101010101" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg341(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"101010110" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg342(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"101010111" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg343(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"101011000" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg344(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"101011001" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg345(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"101011010" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg346(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"101011011" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg347(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"101011100" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg348(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"101011101" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg349(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"101011110" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg350(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"101011111" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg351(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"101100000" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg352(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"101100001" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg353(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"101100010" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg354(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"101100011" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg355(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"101100100" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg356(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"101100101" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg357(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"101100110" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg358(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"101100111" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg359(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"101101000" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg360(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"101101001" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg361(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"101101010" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg362(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"101101011" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg363(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"101101100" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg364(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"101101101" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg365(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"101101110" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg366(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"101101111" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg367(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"101110000" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg368(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"101110001" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg369(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"101110010" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg370(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"101110011" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg371(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"101110100" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg372(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"101110101" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg373(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"101110110" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg374(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"101110111" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg375(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"101111000" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg376(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"101111001" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg377(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"101111010" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg378(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"101111011" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg379(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"101111100" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg380(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"101111101" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg381(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"101111110" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg382(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"101111111" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg383(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"110000000" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg384(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"110000001" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg385(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"110000010" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg386(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"110000011" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg387(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"110000100" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg388(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"110000101" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg389(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"110000110" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg390(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"110000111" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg391(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"110001000" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg392(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"110001001" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg393(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"110001010" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg394(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"110001011" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg395(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"110001100" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg396(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"110001101" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg397(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"110001110" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg398(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"110001111" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg399(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"110010000" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg400(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"110010001" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg401(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"110010010" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg402(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"110010011" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg403(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"110010100" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg404(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"110010101" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg405(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"110010110" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg406(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"110010111" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg407(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"110011000" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg408(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"110011001" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg409(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"110011010" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg410(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"110011011" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg411(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"110011100" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg412(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"110011101" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg413(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"110011110" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg414(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"110011111" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg415(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"110100000" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg416(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"110100001" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg417(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"110100010" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg418(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"110100011" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg419(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"110100100" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg420(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"110100101" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg421(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"110100110" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg422(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"110100111" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg423(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"110101000" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg424(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"110101001" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg425(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"110101010" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg426(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"110101011" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg427(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"110101100" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg428(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"110101101" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg429(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"110101110" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg430(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"110101111" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg431(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"110110000" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg432(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"110110001" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg433(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"110110010" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg434(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"110110011" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg435(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"110110100" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg436(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"110110101" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg437(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"110110110" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg438(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"110110111" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg439(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"110111000" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg440(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"110111001" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg441(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"110111010" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg442(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"110111011" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg443(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"110111100" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg444(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"110111101" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg445(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"110111110" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg446(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"110111111" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg447(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"111000000" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg448(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"111000001" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg449(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"111000010" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg450(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"111000011" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg451(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"111000100" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg452(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"111000101" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg453(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"111000110" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg454(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"111000111" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg455(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"111001000" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg456(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"111001001" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg457(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"111001010" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg458(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"111001011" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg459(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"111001100" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg460(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"111001101" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg461(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"111001110" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg462(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"111001111" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg463(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"111010000" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg464(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"111010001" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg465(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"111010010" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg466(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"111010011" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg467(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"111010100" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg468(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"111010101" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg469(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"111010110" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg470(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"111010111" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg471(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"111011000" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg472(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"111011001" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg473(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"111011010" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg474(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"111011011" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg475(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"111011100" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg476(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"111011101" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg477(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"111011110" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg478(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"111011111" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg479(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"111100000" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg480(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"111100001" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg481(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"111100010" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg482(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"111100011" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg483(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"111100100" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg484(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"111100101" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg485(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"111100110" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg486(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"111100111" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg487(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"111101000" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg488(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"111101001" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg489(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"111101010" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg490(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"111101011" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg491(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"111101100" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg492(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"111101101" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg493(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"111101110" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg494(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"111101111" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg495(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"111110000" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg496(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"111110001" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg497(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"111110010" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg498(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"111110011" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg499(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"111110100" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg500(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"111110101" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg501(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"111110110" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg502(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"111110111" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg503(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"111111000" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg504(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"111111001" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg505(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"111111010" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg506(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"111111011" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg507(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"111111100" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg508(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"111111101" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg509(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"111111110" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg510(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
           when b"111111111" =>      for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop if(S_AXI_WSTRB(byte_index)='1') then        slv_reg511(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);    end if;    end loop;
    when others =>
        slv_reg0<=slv_reg0;     slv_reg1<=slv_reg1;	    slv_reg2<=slv_reg2;	    slv_reg3<=slv_reg3;	
        slv_reg4<=slv_reg4;	    slv_reg5<=slv_reg5;	    slv_reg6<=slv_reg6;	    slv_reg7<=slv_reg7;	
        slv_reg8<=slv_reg8;	    slv_reg9<=slv_reg9;	    slv_reg10<=slv_reg10;	slv_reg11<=slv_reg11;	
        slv_reg12<=slv_reg12;	slv_reg13<=slv_reg13;	slv_reg14<=slv_reg14;	slv_reg15<=slv_reg15;	
        slv_reg16<=slv_reg16;	slv_reg17<=slv_reg17;	slv_reg18<=slv_reg18;	slv_reg19<=slv_reg19;	
        slv_reg20<=slv_reg20;	slv_reg21<=slv_reg21;	slv_reg22<=slv_reg22;	slv_reg23<=slv_reg23;	
        slv_reg24<=slv_reg24;	slv_reg25<=slv_reg25;	slv_reg26<=slv_reg26;	slv_reg27<=slv_reg27;	
        slv_reg28<=slv_reg28;	slv_reg29<=slv_reg29;	slv_reg30<=slv_reg30;	slv_reg31<=slv_reg31;	
        slv_reg32<=slv_reg32;	slv_reg33<=slv_reg33;	slv_reg34<=slv_reg34;	slv_reg35<=slv_reg35;	
        slv_reg36<=slv_reg36;	slv_reg37<=slv_reg37;	slv_reg38<=slv_reg38;	slv_reg39<=slv_reg39;	
        slv_reg40<=slv_reg40;	slv_reg41<=slv_reg41;	slv_reg42<=slv_reg42;	slv_reg43<=slv_reg43;	
        slv_reg44<=slv_reg44;	slv_reg45<=slv_reg45;	slv_reg46<=slv_reg46;	slv_reg47<=slv_reg47;	
        slv_reg48<=slv_reg48;	slv_reg49<=slv_reg49;	slv_reg50<=slv_reg50;	slv_reg51<=slv_reg51;	
        slv_reg52<=slv_reg52;	slv_reg53<=slv_reg53;	slv_reg54<=slv_reg54;	slv_reg55<=slv_reg55;	
        slv_reg56<=slv_reg56;	slv_reg57<=slv_reg57;	slv_reg58<=slv_reg58;	slv_reg59<=slv_reg59;	
        slv_reg60<=slv_reg60;	slv_reg61<=slv_reg61;	slv_reg62<=slv_reg62;	slv_reg63<=slv_reg63;	
        
        slv_reg64<=slv_reg64;	slv_reg65<=slv_reg65;	slv_reg66<=slv_reg66;	slv_reg67<=slv_reg67;	
        slv_reg68<=slv_reg68;	slv_reg69<=slv_reg69;	slv_reg70<=slv_reg70;	slv_reg71<=slv_reg71;	
        slv_reg72<=slv_reg72;	slv_reg73<=slv_reg73;	slv_reg74<=slv_reg74;	slv_reg75<=slv_reg75;	
        slv_reg76<=slv_reg76;	slv_reg77<=slv_reg77;	slv_reg78<=slv_reg78;	slv_reg79<=slv_reg79;	
        slv_reg80<=slv_reg80;	slv_reg81<=slv_reg81;	slv_reg82<=slv_reg82;	slv_reg83<=slv_reg83;	
        slv_reg84<=slv_reg84;	slv_reg85<=slv_reg85;	slv_reg86<=slv_reg86;	slv_reg87<=slv_reg87;	
        slv_reg88<=slv_reg88;	slv_reg89<=slv_reg89;	slv_reg90<=slv_reg90;	slv_reg91<=slv_reg91;	
        slv_reg92<=slv_reg92;	slv_reg93<=slv_reg93;	slv_reg94<=slv_reg94;	slv_reg95<=slv_reg95;	
        slv_reg96<=slv_reg96;	slv_reg97<=slv_reg97;	slv_reg98<=slv_reg98;	slv_reg99<=slv_reg99;	
        slv_reg100<=slv_reg100;	slv_reg101<=slv_reg101;	slv_reg102<=slv_reg102;	slv_reg103<=slv_reg103;	
        slv_reg104<=slv_reg104;	slv_reg105<=slv_reg105;	slv_reg106<=slv_reg106;	slv_reg107<=slv_reg107;	
        slv_reg108<=slv_reg108;	slv_reg109<=slv_reg109;	slv_reg110<=slv_reg110;	slv_reg111<=slv_reg111;	
        slv_reg112<=slv_reg112;	slv_reg113<=slv_reg113;	slv_reg114<=slv_reg114;	slv_reg115<=slv_reg115;	
        slv_reg116<=slv_reg116;	slv_reg117<=slv_reg117;	slv_reg118<=slv_reg118;	slv_reg119<=slv_reg119;	
        slv_reg120<=slv_reg120;	slv_reg121<=slv_reg121;	slv_reg122<=slv_reg122;	slv_reg123<=slv_reg123;	
        slv_reg124<=slv_reg124;	slv_reg125<=slv_reg125;	slv_reg126<=slv_reg126;	slv_reg127<=slv_reg127;
        	
        slv_reg128<=slv_reg128;	slv_reg129<=slv_reg129;	slv_reg130<=slv_reg130;	slv_reg131<=slv_reg131;	
        slv_reg132<=slv_reg132;	slv_reg133<=slv_reg133;	slv_reg134<=slv_reg134;	slv_reg135<=slv_reg135;	
        slv_reg136<=slv_reg136;	slv_reg137<=slv_reg137;	slv_reg138<=slv_reg138;	slv_reg139<=slv_reg139;	
        slv_reg140<=slv_reg140;	slv_reg141<=slv_reg141;	slv_reg142<=slv_reg142;	slv_reg143<=slv_reg143;	
        slv_reg144<=slv_reg144;	slv_reg145<=slv_reg145;	slv_reg146<=slv_reg146;	slv_reg147<=slv_reg147;	
        slv_reg148<=slv_reg148;	slv_reg149<=slv_reg149;	slv_reg150<=slv_reg150;	slv_reg151<=slv_reg151;	
        slv_reg152<=slv_reg152;	slv_reg153<=slv_reg153;	slv_reg154<=slv_reg154;	slv_reg155<=slv_reg155;	
        slv_reg156<=slv_reg156;	slv_reg157<=slv_reg157;	slv_reg158<=slv_reg158;	slv_reg159<=slv_reg159;	
        slv_reg160<=slv_reg160;	slv_reg161<=slv_reg161;	slv_reg162<=slv_reg162;	slv_reg163<=slv_reg163;	
        slv_reg164<=slv_reg164;	slv_reg165<=slv_reg165;	slv_reg166<=slv_reg166;	slv_reg167<=slv_reg167;	
        slv_reg168<=slv_reg168;	slv_reg169<=slv_reg169;	slv_reg170<=slv_reg170;	slv_reg171<=slv_reg171;
        slv_reg172<=slv_reg172;	slv_reg173<=slv_reg173;	slv_reg174<=slv_reg174;	slv_reg175<=slv_reg175;	
        slv_reg176<=slv_reg176;	slv_reg177<=slv_reg177;	slv_reg178<=slv_reg178;	slv_reg179<=slv_reg179;	
        slv_reg180<=slv_reg180;	slv_reg181<=slv_reg181;	slv_reg182<=slv_reg182;	slv_reg183<=slv_reg183;	
        slv_reg184<=slv_reg184;	slv_reg185<=slv_reg185;	slv_reg186<=slv_reg186;	slv_reg187<=slv_reg187;	
        slv_reg188<=slv_reg188;	slv_reg189<=slv_reg189;	slv_reg190<=slv_reg190;	slv_reg191<=slv_reg191;
              
        slv_reg192<=slv_reg192;	slv_reg193<=slv_reg193;	slv_reg194<=slv_reg194;	slv_reg195<=slv_reg195;	
        slv_reg196<=slv_reg196;	slv_reg197<=slv_reg197;	slv_reg198<=slv_reg198;	slv_reg199<=slv_reg199;	
        slv_reg200<=slv_reg200;	slv_reg201<=slv_reg201;	slv_reg202<=slv_reg202;	slv_reg203<=slv_reg203;	
        slv_reg204<=slv_reg204;	slv_reg205<=slv_reg205;	slv_reg206<=slv_reg206;	slv_reg207<=slv_reg207;	
        slv_reg208<=slv_reg208;	slv_reg209<=slv_reg209;	slv_reg210<=slv_reg210;	slv_reg211<=slv_reg211;	
        slv_reg212<=slv_reg212;	slv_reg213<=slv_reg213;	slv_reg214<=slv_reg214;	slv_reg215<=slv_reg215;	
        slv_reg216<=slv_reg216;	slv_reg217<=slv_reg217;	slv_reg218<=slv_reg218;	slv_reg219<=slv_reg219;	
        slv_reg220<=slv_reg220;	slv_reg221<=slv_reg221;	slv_reg222<=slv_reg222;	slv_reg223<=slv_reg223;	
        slv_reg224<=slv_reg224;	slv_reg225<=slv_reg225;	slv_reg226<=slv_reg226;	slv_reg227<=slv_reg227;	
        slv_reg228<=slv_reg228;	slv_reg229<=slv_reg229;	slv_reg230<=slv_reg230;	slv_reg231<=slv_reg231;	
        slv_reg232<=slv_reg232;	slv_reg233<=slv_reg233;	slv_reg234<=slv_reg234;	slv_reg235<=slv_reg235;	
        slv_reg236<=slv_reg236;	slv_reg237<=slv_reg237;	slv_reg238<=slv_reg238;	slv_reg239<=slv_reg239;	
        slv_reg240<=slv_reg240;	slv_reg241<=slv_reg241;	slv_reg242<=slv_reg242;	slv_reg243<=slv_reg243;	
        slv_reg244<=slv_reg244;	slv_reg245<=slv_reg245;	slv_reg246<=slv_reg246;	slv_reg247<=slv_reg247;	
        slv_reg248<=slv_reg248;	slv_reg249<=slv_reg249;	slv_reg250<=slv_reg250;	slv_reg251<=slv_reg251;	
        slv_reg252<=slv_reg252;	slv_reg253<=slv_reg253;	slv_reg254<=slv_reg254;	slv_reg255<=slv_reg255;
        	
        slv_reg256<=slv_reg256;	slv_reg257<=slv_reg257;	slv_reg258<=slv_reg258;	slv_reg259<=slv_reg259;	
        slv_reg260<=slv_reg260;	slv_reg261<=slv_reg261;	slv_reg262<=slv_reg262;	slv_reg263<=slv_reg263;	
        slv_reg264<=slv_reg264;	slv_reg265<=slv_reg265;	slv_reg266<=slv_reg266;	slv_reg267<=slv_reg267;	
        slv_reg268<=slv_reg268;	slv_reg269<=slv_reg269;	slv_reg270<=slv_reg270;	slv_reg271<=slv_reg271;	
        slv_reg272<=slv_reg272;	slv_reg273<=slv_reg273;	slv_reg274<=slv_reg274;	slv_reg275<=slv_reg275;	
        slv_reg276<=slv_reg276;	slv_reg277<=slv_reg277;	slv_reg278<=slv_reg278;	slv_reg279<=slv_reg279;	
        slv_reg280<=slv_reg280;	slv_reg281<=slv_reg281;	slv_reg282<=slv_reg282;	slv_reg283<=slv_reg283;	
        slv_reg284<=slv_reg284;	slv_reg285<=slv_reg285;	slv_reg286<=slv_reg286;	slv_reg287<=slv_reg287;	
        slv_reg288<=slv_reg288;	slv_reg289<=slv_reg289;	slv_reg290<=slv_reg290;	slv_reg291<=slv_reg291;
        slv_reg292<=slv_reg292;	slv_reg293<=slv_reg293;	slv_reg294<=slv_reg294;	slv_reg295<=slv_reg295;	
        slv_reg296<=slv_reg296;	slv_reg297<=slv_reg297;	slv_reg298<=slv_reg298;	slv_reg299<=slv_reg299;	
        slv_reg300<=slv_reg300;	slv_reg301<=slv_reg301;	slv_reg302<=slv_reg302;	slv_reg303<=slv_reg303;	
        slv_reg304<=slv_reg304;	slv_reg305<=slv_reg305;	slv_reg306<=slv_reg306;	slv_reg307<=slv_reg307;	
        slv_reg308<=slv_reg308;	slv_reg309<=slv_reg309;	slv_reg310<=slv_reg310;	slv_reg311<=slv_reg311;	
        slv_reg312<=slv_reg312;	slv_reg313<=slv_reg313;	slv_reg314<=slv_reg314;	slv_reg315<=slv_reg315;	
        slv_reg316<=slv_reg316;	slv_reg317<=slv_reg317;	slv_reg318<=slv_reg318;	slv_reg319<=slv_reg319;
        	
        slv_reg320<=slv_reg320;	slv_reg321<=slv_reg321;	slv_reg322<=slv_reg322;	slv_reg323<=slv_reg323;	
        slv_reg324<=slv_reg324;	slv_reg325<=slv_reg325;	slv_reg326<=slv_reg326;	slv_reg327<=slv_reg327;	
        slv_reg328<=slv_reg328;	slv_reg329<=slv_reg329;	slv_reg330<=slv_reg330;	slv_reg331<=slv_reg331;	
        slv_reg332<=slv_reg332;	slv_reg333<=slv_reg333;	slv_reg334<=slv_reg334;	slv_reg335<=slv_reg335;	
        slv_reg336<=slv_reg336;	slv_reg337<=slv_reg337;	slv_reg338<=slv_reg338;	slv_reg339<=slv_reg339;	
        slv_reg340<=slv_reg340;	slv_reg341<=slv_reg341;	slv_reg342<=slv_reg342;	slv_reg343<=slv_reg343;	
        slv_reg344<=slv_reg344;	slv_reg345<=slv_reg345;	slv_reg346<=slv_reg346;	slv_reg347<=slv_reg347;	
        slv_reg348<=slv_reg348;	slv_reg349<=slv_reg349;	slv_reg350<=slv_reg350;	slv_reg351<=slv_reg351;	
        slv_reg352<=slv_reg352;	slv_reg353<=slv_reg353;	slv_reg354<=slv_reg354;	slv_reg355<=slv_reg355;	
        slv_reg356<=slv_reg356;	slv_reg357<=slv_reg357;	slv_reg358<=slv_reg358;	slv_reg359<=slv_reg359;	
        slv_reg360<=slv_reg360;	slv_reg361<=slv_reg361;	slv_reg362<=slv_reg362;	slv_reg363<=slv_reg363;	
        slv_reg364<=slv_reg364;	slv_reg365<=slv_reg365;	slv_reg366<=slv_reg366;	slv_reg367<=slv_reg367;	
        slv_reg368<=slv_reg368;	slv_reg369<=slv_reg369;	slv_reg370<=slv_reg370;	slv_reg371<=slv_reg371;	
        slv_reg372<=slv_reg372;	slv_reg373<=slv_reg373;	slv_reg374<=slv_reg374;	slv_reg375<=slv_reg375;	
        slv_reg376<=slv_reg376;	slv_reg377<=slv_reg377;	slv_reg378<=slv_reg378;	slv_reg379<=slv_reg379;	
        slv_reg380<=slv_reg380;	slv_reg381<=slv_reg381;	slv_reg382<=slv_reg382;	slv_reg383<=slv_reg383;
        	
        slv_reg384<=slv_reg384;	slv_reg385<=slv_reg385;	slv_reg386<=slv_reg386;	slv_reg387<=slv_reg387;	
        slv_reg388<=slv_reg388;	slv_reg389<=slv_reg389;	slv_reg390<=slv_reg390;	slv_reg391<=slv_reg391;	
        slv_reg392<=slv_reg392;	slv_reg393<=slv_reg393;	slv_reg394<=slv_reg394;	slv_reg395<=slv_reg395;	
        slv_reg396<=slv_reg396;	slv_reg397<=slv_reg397;	slv_reg398<=slv_reg398;	slv_reg399<=slv_reg399;	
        slv_reg400<=slv_reg400;	slv_reg401<=slv_reg401;	slv_reg402<=slv_reg402;	slv_reg403<=slv_reg403;	
        slv_reg404<=slv_reg404;	slv_reg405<=slv_reg405;	slv_reg406<=slv_reg406;	slv_reg407<=slv_reg407;
        slv_reg408<=slv_reg408;	slv_reg409<=slv_reg409;	slv_reg410<=slv_reg410;	slv_reg411<=slv_reg411;	
        slv_reg412<=slv_reg412;	slv_reg413<=slv_reg413;	slv_reg414<=slv_reg414;	slv_reg415<=slv_reg415;	
        slv_reg416<=slv_reg416;	slv_reg417<=slv_reg417;	slv_reg418<=slv_reg418;	slv_reg419<=slv_reg419;	
        slv_reg420<=slv_reg420;	slv_reg421<=slv_reg421;	slv_reg422<=slv_reg422;	slv_reg423<=slv_reg423;	
        slv_reg424<=slv_reg424;	slv_reg425<=slv_reg425;	slv_reg426<=slv_reg426;	slv_reg427<=slv_reg427;	
        slv_reg428<=slv_reg428;	slv_reg429<=slv_reg429;	slv_reg430<=slv_reg430;	slv_reg431<=slv_reg431;	
        slv_reg432<=slv_reg432;	slv_reg433<=slv_reg433;	slv_reg434<=slv_reg434;	slv_reg435<=slv_reg435;	
        slv_reg436<=slv_reg436;	slv_reg437<=slv_reg437;	slv_reg438<=slv_reg438;	slv_reg439<=slv_reg439;	
        slv_reg440<=slv_reg440;	slv_reg441<=slv_reg441;	slv_reg442<=slv_reg442;	slv_reg443<=slv_reg443;	
        slv_reg444<=slv_reg444;	slv_reg445<=slv_reg445;	slv_reg446<=slv_reg446;	slv_reg447<=slv_reg447;
        	
        slv_reg448<=slv_reg448;	slv_reg449<=slv_reg449;	slv_reg450<=slv_reg450;	slv_reg451<=slv_reg451;	
        slv_reg452<=slv_reg452;	slv_reg453<=slv_reg453;	slv_reg454<=slv_reg454;	slv_reg455<=slv_reg455;	
        slv_reg456<=slv_reg456;	slv_reg457<=slv_reg457;	slv_reg458<=slv_reg458;	slv_reg459<=slv_reg459;	
        slv_reg460<=slv_reg460;	slv_reg461<=slv_reg461;	slv_reg462<=slv_reg462;	slv_reg463<=slv_reg463;	
        slv_reg464<=slv_reg464;	slv_reg465<=slv_reg465;	slv_reg466<=slv_reg466;	slv_reg467<=slv_reg467;	
        slv_reg468<=slv_reg468;	slv_reg469<=slv_reg469;	slv_reg470<=slv_reg470;	slv_reg471<=slv_reg471;	
        slv_reg472<=slv_reg472;	slv_reg473<=slv_reg473;	slv_reg474<=slv_reg474;	slv_reg475<=slv_reg475;	
        slv_reg476<=slv_reg476;	slv_reg477<=slv_reg477;	slv_reg478<=slv_reg478;	slv_reg479<=slv_reg479;	
        slv_reg480<=slv_reg480;	slv_reg481<=slv_reg481;	slv_reg482<=slv_reg482;	slv_reg483<=slv_reg483;	
        slv_reg484<=slv_reg484;	slv_reg485<=slv_reg485;	slv_reg486<=slv_reg486;	slv_reg487<=slv_reg487;	
        slv_reg488<=slv_reg488;	slv_reg489<=slv_reg489;	slv_reg490<=slv_reg490;	slv_reg491<=slv_reg491;	
        slv_reg492<=slv_reg492;	slv_reg493<=slv_reg493;	slv_reg494<=slv_reg494;	slv_reg495<=slv_reg495;	
        slv_reg496<=slv_reg496;	slv_reg497<=slv_reg497;	slv_reg498<=slv_reg498;	slv_reg499<=slv_reg499;	
        slv_reg500<=slv_reg500;	slv_reg501<=slv_reg501;	slv_reg502<=slv_reg502;	slv_reg503<=slv_reg503;	
        slv_reg504<=slv_reg504;	slv_reg505<=slv_reg505;	slv_reg506<=slv_reg506;	slv_reg507<=slv_reg507;	
        slv_reg508<=slv_reg508;	slv_reg509<=slv_reg509;	slv_reg510<=slv_reg510;	slv_reg511<=slv_reg511;
    end case;
    end if;    end if;    end if;       end process; 

	process (S_AXI_ACLK)
	begin
	  if rising_edge(S_AXI_ACLK) then 
	    if S_AXI_ARESETN = '0' then
	      axi_bvalid <='0';
	      axi_bresp  <="00"; --need to work more on the responses
	    else
	      if (axi_awready = '1' and S_AXI_AWVALID = '1' and axi_wready = '1' and S_AXI_WVALID = '1' and axi_bvalid = '0'  ) then
	        axi_bvalid<='1';
	        axi_bresp <="00"; 
	      elsif (S_AXI_BREADY = '1' and axi_bvalid = '1') then   --check if bready is asserted while bvalid is high)
	        axi_bvalid<='0';                                 -- (there is a possibility that bready is always asserted high)
	      end if;
	    end if;
	  end if;                   
	end process; 

	process (S_AXI_ACLK)
	begin
	  if rising_edge(S_AXI_ACLK) then 
	    if S_AXI_ARESETN = '0' then
	      axi_arready<='0';
	      axi_araddr <=(others => '1');
	    else
	      if (axi_arready = '0' and S_AXI_ARVALID = '1') then
	        -- indicates that the slave has acceped the valid read address
	        axi_arready <= '1';
	        -- Read Address latching 
	        axi_araddr  <= S_AXI_ARADDR;           
	      else
	        axi_arready <= '0';
	      end if;
	    end if;
	  end if;                   
	end process; 

	process (S_AXI_ACLK)
	begin
	  if rising_edge(S_AXI_ACLK) then
	    if S_AXI_ARESETN = '0' then
	      axi_rvalid <= '0';
	      axi_rresp  <= "00";
	    else
	      if (axi_arready = '1' and S_AXI_ARVALID = '1' and axi_rvalid = '0') then
	        axi_rvalid <= '1';
	        axi_rresp  <= "00"; -- 'OKAY' response
	      elsif (axi_rvalid = '1' and S_AXI_RREADY = '1') then
	        axi_rvalid <= '0';
	      end if;            
	    end if;
	  end if;
	end process;
	slv_reg_rden <= axi_arready and S_AXI_ARVALID and (not axi_rvalid) ;
    
    -- Output register or memory read data
        process( S_AXI_ACLK ) is
        begin
          if (rising_edge (S_AXI_ACLK)) then
            if ( S_AXI_ARESETN = '0' ) then
              axi_rdata  <= (others => '0');
            else
              if (slv_reg_rden = '1') then
                axi_rdata <= reg_data_out;     -- register read data
              end if;   
            end if;
          end if;
        end process;
    
    






end arch_imp;
